// Generator : SpinalHDL dev    git head : 93c1ed9a2922adbb6c8bf1ba3a8a0a652c1b8bbf
// Component : VexiiRiscv
// Git hash  : 74c61a50ae672f9f203188a850dc54e1ca50ca08

`timescale 1ns/1ps

module VexiiRiscv (
  input  wire [63:0]   PrivilegedPlugin_logic_rdtime,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_timer /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_software /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_external /* verilator public */ ,
  output wire          LsuL1WishbonePlugin_logic_bus_CYC,
  output wire          LsuL1WishbonePlugin_logic_bus_STB,
  input  wire          LsuL1WishbonePlugin_logic_bus_ACK,
  output wire          LsuL1WishbonePlugin_logic_bus_WE,
  output wire [26:0]   LsuL1WishbonePlugin_logic_bus_ADR,
  input  wire [255:0]  LsuL1WishbonePlugin_logic_bus_DAT_MISO,
  output wire [255:0]  LsuL1WishbonePlugin_logic_bus_DAT_MOSI,
  output wire [31:0]   LsuL1WishbonePlugin_logic_bus_SEL,
  input  wire          LsuL1WishbonePlugin_logic_bus_ERR,
  output wire [2:0]    LsuL1WishbonePlugin_logic_bus_CTI,
  output wire [1:0]    LsuL1WishbonePlugin_logic_bus_BTE,
  output reg           FetchL1WishbonePlugin_logic_bus_CYC,
  output reg           FetchL1WishbonePlugin_logic_bus_STB,
  input  wire          FetchL1WishbonePlugin_logic_bus_ACK,
  output wire          FetchL1WishbonePlugin_logic_bus_WE,
  output wire [26:0]   FetchL1WishbonePlugin_logic_bus_ADR,
  input  wire [255:0]  FetchL1WishbonePlugin_logic_bus_DAT_MISO,
  output wire [255:0]  FetchL1WishbonePlugin_logic_bus_DAT_MOSI,
  output wire [31:0]   FetchL1WishbonePlugin_logic_bus_SEL,
  input  wire          FetchL1WishbonePlugin_logic_bus_ERR,
  output wire [2:0]    FetchL1WishbonePlugin_logic_bus_CTI,
  output wire [1:0]    FetchL1WishbonePlugin_logic_bus_BTE,
  output wire          LsuCachelessWishbonePlugin_logic_bridge_down_CYC,
  output wire          LsuCachelessWishbonePlugin_logic_bridge_down_STB,
  input  wire          LsuCachelessWishbonePlugin_logic_bridge_down_ACK,
  output wire          LsuCachelessWishbonePlugin_logic_bridge_down_WE,
  output wire [28:0]   LsuCachelessWishbonePlugin_logic_bridge_down_ADR,
  input  wire [63:0]   LsuCachelessWishbonePlugin_logic_bridge_down_DAT_MISO,
  output wire [63:0]   LsuCachelessWishbonePlugin_logic_bridge_down_DAT_MOSI,
  output wire [7:0]    LsuCachelessWishbonePlugin_logic_bridge_down_SEL,
  input  wire          LsuCachelessWishbonePlugin_logic_bridge_down_ERR,
  output wire [2:0]    LsuCachelessWishbonePlugin_logic_bridge_down_CTI,
  output wire [1:0]    LsuCachelessWishbonePlugin_logic_bridge_down_BTE,
  input  wire          clk,
  input  wire          reset
);
  localparam FloatMode_ZERO = 2'd0;
  localparam FloatMode_INF = 2'd1;
  localparam FloatMode_NAN = 2'd2;
  localparam FloatMode_NORMAL = 2'd3;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;
  localparam FpuFormat_FpuCmpPlugin_logic_f32_1 = 1'd0;
  localparam FpuFormat_FpuCmpPlugin_logic_f64_1 = 1'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_ZERO = 2'd3;
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam FpuCmpFloatOp_MIN_MAX = 1'd0;
  localparam FpuCmpFloatOp_SGNJ = 1'd1;
  localparam EnvPluginOp_ECALL = 3'd0;
  localparam EnvPluginOp_EBREAK = 3'd1;
  localparam EnvPluginOp_PRIV_RET = 3'd2;
  localparam EnvPluginOp_FENCE_I = 3'd3;
  localparam EnvPluginOp_SFENCE_VMA = 3'd4;
  localparam EnvPluginOp_WFI = 3'd5;
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;
  localparam LsuPlugin_logic_flusher_IDLE = 2'd0;
  localparam LsuPlugin_logic_flusher_SB_DRAIN = 2'd1;
  localparam LsuPlugin_logic_flusher_CMD = 2'd2;
  localparam LsuPlugin_logic_flusher_COMPLETION = 2'd3;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RESET = 4'd0;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RUNNING = 4'd1;
  localparam TrapPlugin_logic_harts_0_trap_fsm_COMPUTE = 4'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC = 4'd3;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL = 4'd4;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC = 4'd5;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY = 4'd6;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC = 4'd7;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY = 4'd8;
  localparam TrapPlugin_logic_harts_0_trap_fsm_JUMP = 4'd9;
  localparam TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH = 4'd10;
  localparam TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH = 4'd11;
  localparam CsrAccessPlugin_logic_fsm_IDLE = 2'd0;
  localparam CsrAccessPlugin_logic_fsm_READ = 2'd1;
  localparam CsrAccessPlugin_logic_fsm_WRITE = 2'd2;
  localparam CsrAccessPlugin_logic_fsm_COMPLETION = 2'd3;

  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_ready;
  reg                 FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid;
  reg        [51:0]   FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data;
  wire                FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_valid;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_payload_data;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_valid;
  reg                 early0_DivPlugin_logic_processing_div_io_cmd_payload_normalized;
  reg        [4:0]    early0_DivPlugin_logic_processing_div_io_cmd_payload_iterations;
  reg                 LsuPlugin_logic_flusher_arbiter_io_output_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_ready;
  wire                FpuSqrtPlugin_logic_sqrt_io_input_valid;
  wire       [53:0]   FpuSqrtPlugin_logic_sqrt_io_input_payload_a;
  reg                 integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid;
  reg        [4:0]    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address;
  reg        [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data;
  reg                 float_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid;
  reg        [4:0]    float_RegFilePlugin_logic_regfile_fpga_io_writes_0_address;
  reg        [63:0]   float_RegFilePlugin_logic_regfile_fpga_io_writes_0_data;
  wire       [30:0]   BtbPlugin_logic_ras_mem_stack_spinal_port0;
  reg        [255:0]  LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [255:0]  LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [2:0]    LsuL1Plugin_logic_shared_mem_spinal_port1;
  reg        [255:0]  LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  reg        [51:0]   PrefetcherRptPlugin_logic_storage_ram_spinal_port0;
  reg        [255:0]  FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [255:0]  FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [0:0]    FetchL1Plugin_logic_plru_mem_spinal_port1;
  reg        [7:0]    GSharePlugin_logic_mem_banks_0_spinal_port1;
  reg        [93:0]   BtbPlugin_logic_mem_spinal_port1;
  reg        [109:0]  LsuPlugin_logic_storeBuffer_ops_mem_spinal_port0;
  reg        [31:0]   CsrRamPlugin_logic_mem_spinal_port1;
  wire                PrefetcherRptPlugin_logic_order_fifo_io_push_ready;
  wire                PrefetcherRptPlugin_logic_order_fifo_io_pop_valid;
  wire       [31:0]   PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_address;
  wire                PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_stride;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_fifo_io_occupancy;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_fifo_io_availability;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_0_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_1_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_valid;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_last;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_write;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_id;
  wire       [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_address;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_chosen;
  wire       [1:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_chosenOH;
  wire                FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_ready;
  wire                FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_ready;
  wire                FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_valid;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_payload_data;
  wire       [0:0]    FpuUnpackerPlugin_logic_unpacker_arbiter_io_chosen;
  wire       [1:0]    FpuUnpackerPlugin_logic_unpacker_arbiter_io_chosenOH;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_ready;
  wire                early0_DivPlugin_logic_processing_div_io_rsp_valid;
  wire       [63:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_result;
  wire       [63:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_remain;
  wire                LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_flusher_arbiter_io_output_valid;
  wire       [0:0]    LsuPlugin_logic_flusher_arbiter_io_chosenOH;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_3_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosen;
  wire       [3:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosenOH;
  wire                streamArbiter_5_io_inputs_0_ready;
  wire                streamArbiter_5_io_inputs_1_ready;
  wire                streamArbiter_5_io_output_valid;
  wire       [31:0]   streamArbiter_5_io_output_payload_pcOnLastSlice;
  wire       [31:0]   streamArbiter_5_io_output_payload_pcTarget;
  wire                streamArbiter_5_io_output_payload_taken;
  wire                streamArbiter_5_io_output_payload_isBranch;
  wire                streamArbiter_5_io_output_payload_isPush;
  wire                streamArbiter_5_io_output_payload_isPop;
  wire                streamArbiter_5_io_output_payload_wasWrong;
  wire                streamArbiter_5_io_output_payload_badPredictedTarget;
  wire       [11:0]   streamArbiter_5_io_output_payload_history;
  wire       [15:0]   streamArbiter_5_io_output_payload_uopId;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire       [0:0]    streamArbiter_5_io_chosen;
  wire       [1:0]    streamArbiter_5_io_chosenOH;
  wire                FpuSqrtPlugin_logic_sqrt_io_input_ready;
  wire                FpuSqrtPlugin_logic_sqrt_io_output_valid;
  wire       [52:0]   FpuSqrtPlugin_logic_sqrt_io_output_payload_result;
  wire       [56:0]   FpuSqrtPlugin_logic_sqrt_io_output_payload_remain;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
  wire       [63:0]   float_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [63:0]   float_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [63:0]   float_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early0_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_1_mem_port_1;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_mem_port;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_refill_free_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_refill_free_2;
  reg        [25:0]   _zz_LsuL1Plugin_logic_refill_read_cmdAddress;
  reg        [31:0]   _zz_LsuL1Plugin_logic_refill_read_rspAddress;
  reg                 _zz_LsuL1Plugin_logic_refill_read_dirty;
  reg        [0:0]    _zz_LsuL1Plugin_logic_refill_read_way;
  wire       [1:0]    _zz_LsuL1Plugin_logic_writeback_free_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_writeback_free_2;
  reg        [31:0]   _zz_LsuL1Plugin_logic_writeback_read_address;
  reg        [0:0]    _zz_LsuL1Plugin_logic_writeback_read_way;
  reg        [255:0]  _zz_LsuL1Plugin_logic_writeback_read_readedData;
  wire       [1:0]    _zz_LsuL1Plugin_logic_writeback_victimBuffer_port;
  reg        [31:0]   _zz_LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  reg        [63:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [1:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1;
  reg        [63:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [0:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite;
  reg        [1:0]    _zz_59;
  wire       [1:0]    _zz_60;
  reg        [1:0]    _zz_61;
  wire       [2:0]    _zz_62;
  wire       [1:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty;
  reg        [19:0]   _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
  reg        [19:0]   _zz_LsuL1Plugin_logic_writeback_push_payload_address;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1;
  wire       [2:0]    _zz_PrefetcherRptPlugin_logic_counter;
  wire       [2:0]    _zz_PrefetcherRptPlugin_logic_counter_1;
  wire       [0:0]    _zz_PrefetcherRptPlugin_logic_counter_2;
  wire       [3:0]    _zz_PrefetcherRptPlugin_logic_pip2_node_0_MUL;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_1;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_2;
  wire       [51:0]   _zz_PrefetcherRptPlugin_logic_storage_ram_port;
  wire       [31:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_late0_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_late0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_late0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_late0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_late0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_late0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_late0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_late0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early1_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_early1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_early1_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_early1_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_early1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_early1_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_early1_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_early1_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_late1_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_late1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_late1_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_late1_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_late1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_late1_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_late1_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_late1_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_1_mem_port_1;
  wire                _zz_when;
  wire       [1:0]    _zz_when_1;
  wire       [1:0]    _zz_when_2;
  wire       [0:0]    _zz_FetchL1Plugin_logic_bus_cmd_payload_io;
  wire       [0:0]    _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts;
  wire       [0:0]    _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_1;
  wire       [0:0]    _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_2;
  wire       [0:0]    _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_3;
  reg        [0:0]    _zz_FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  reg        [31:0]   _zz_FetchL1Plugin_logic_refill_onRsp_address;
  reg        [63:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [1:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1;
  reg        [63:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [1:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_dataAccessFault;
  wire       [0:0]    _zz_FetchL1Plugin_logic_plru_write_payload_data_0;
  wire       [7:0]    _zz_GSharePlugin_logic_mem_banks_0_port;
  wire       [1:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1;
  wire       [11:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_4;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4;
  wire       [30:0]   _zz_BtbPlugin_logic_ras_mem_stack_port;
  wire       [93:0]   _zz_BtbPlugin_logic_mem_port;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_1_pc;
  wire       [0:0]    _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire       [25:0]   _zz_FetchL1WishbonePlugin_logic_bus_ADR;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [11:0]   _zz__zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [31:0]   _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3;
  wire       [11:0]   _zz__zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1;
  wire       [31:0]   _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent_1;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent_1;
  wire       [51:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa;
  reg        [1:0]    _zz_63;
  wire       [1:0]    _zz_64;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_2;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_3;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_4;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_2;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_3;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_4;
  wire       [12:0]   _zz__zz_when_AFix_l1168;
  wire       [12:0]   _zz__zz_when_AFix_l1168_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_1;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_2;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_1;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_2;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_3;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_4;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_1;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_2;
  wire       [104:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_3;
  wire       [105:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_4;
  wire       [107:0]  _zz__zz_when_Utils_l1585_13;
  wire       [107:0]  _zz__zz_when_Utils_l1585_12;
  wire       [107:0]  _zz__zz_when_Utils_l1585_11;
  wire       [107:0]  _zz__zz_when_Utils_l1585_10;
  wire       [107:0]  _zz__zz_when_Utils_l1585_9;
  wire       [107:0]  _zz__zz_when_Utils_l1585_8;
  wire       [107:0]  _zz__zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_2;
  wire       [0:0]    _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_3;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_1;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_2;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_1;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_2;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_3;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_4;
  wire       [0:0]    _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_5;
  wire       [108:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa;
  wire       [108:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_1;
  wire       [108:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_2;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_3;
  wire       [106:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_4;
  wire       [108:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_5;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_6;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1;
  wire       [98:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4;
  wire       [87:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7;
  wire       [76:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10;
  wire       [65:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13;
  wire       [54:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16;
  wire       [43:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19;
  wire       [32:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22;
  wire       [21:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24;
  wire       [0:0]    _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25;
  wire       [10:0]   _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_2;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_2;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_2;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_2;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105_1;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106;
  wire                _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_2;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_3;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_4;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_5;
  wire       [7:0]    _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_6;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_7;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_8;
  wire       [108:0]  _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent_1;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_exponent;
  wire       [11:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_exponent;
  wire       [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy;
  wire       [0:0]    _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1;
  wire       [42:0]   _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3;
  wire       [0:0]    _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4;
  wire       [31:0]   _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6;
  wire       [0:0]    _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7;
  wire       [20:0]   _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9;
  wire       [0:0]    _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10;
  wire       [9:0]    _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127;
  wire                _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128;
  wire       [53:0]   _zz_execute_ctrl2_down_MUL_SRC1_lane0;
  wire       [32:0]   _zz_execute_ctrl2_down_MUL_SRC1_lane0_1;
  wire       [53:0]   _zz_execute_ctrl2_down_MUL_SRC2_lane0;
  wire       [32:0]   _zz_execute_ctrl2_down_MUL_SRC2_lane0_1;
  wire       [56:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3;
  wire       [56:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3;
  wire       [39:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3;
  wire       [39:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3;
  wire       [22:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3;
  wire       [22:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [20:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3;
  wire       [5:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17;
  wire       [63:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17;
  wire       [46:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17;
  wire       [5:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18;
  wire       [31:0]   _zz_early0_DivPlugin_logic_processing_selected;
  wire       [31:0]   _zz_early0_DivPlugin_logic_processing_selected_1;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3;
  wire       [3:0]    _zz_early0_EnvPlugin_logic_trapPort_payload_code;
  wire       [20:0]   _zz_early0_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early0_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early0_BranchPlugin_pcCalc_target_b_2;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [2:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [1:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1;
  wire       [20:0]   _zz_early1_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early1_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early1_BranchPlugin_pcCalc_target_b_2;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire       [2:0]    _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire       [1:0]    _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1;
  reg        [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  wire       [1:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1;
  reg        [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2;
  wire       [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_15;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_16;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_17;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_18;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_19;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_20;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_21;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_22;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_24;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_5;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_6;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_15;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_2;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_15;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_16;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_17;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_18;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_19;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_5;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_6;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_11;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26;
  wire       [11:0]   _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
  wire       [5:0]    _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1;
  reg        [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29;
  wire       [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30;
  wire       [6:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_37;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_38;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_39;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_40;
  wire       [1:0]    _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26;
  wire       [11:0]   _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
  wire       [5:0]    _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1;
  reg        [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29;
  wire       [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30;
  wire       [6:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_37;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_38;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_39;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_40;
  wire       [1:0]    _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  wire       [9:0]    _zz_decode_ctrls_0_up_Decode_DOP_ID_1;
  wire       [0:0]    _zz_decode_ctrls_0_up_Decode_DOP_ID_1_1;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice;
  wire       [5:0]    _zz_LsuPlugin_logic_storeBuffer_ops_popPtr;
  wire       [0:0]    _zz_LsuPlugin_logic_storeBuffer_ops_popPtr_1;
  wire       [4:0]    _zz_LsuPlugin_logic_storeBuffer_ops_mem_port;
  wire       [4:0]    _zz__zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1;
  wire       [5:0]    _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr;
  wire       [0:0]    _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr_1;
  wire                _zz_when_3;
  wire                _zz_when_4;
  wire                _zz_when_5;
  wire                _zz_when_6;
  wire                _zz_when_7;
  wire                _zz_when_8;
  wire                _zz_when_9;
  wire                _zz_when_10;
  wire       [4:0]    _zz_LsuPlugin_logic_storeBuffer_ops_mem_port_1;
  wire       [109:0]  _zz_LsuPlugin_logic_storeBuffer_ops_mem_port_2;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_ls_storeId;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_ls_storeId_1;
  wire       [12:0]   _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_5;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_7;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5;
  wire                _zz_LsuPlugin_logic_onCtrl_wb_hits;
  wire                _zz_LsuPlugin_logic_onCtrl_wb_hits_1;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_wb_hits_2;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_wb_hits_3;
  wire       [2:0]    _zz_LsuPlugin_logic_trapPort_payload_code;
  wire                _zz_execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire                _zz_execute_ctrl4_down_LsuL1_ABORD_lane0_1;
  wire                _zz_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0;
  wire       [5:0]    _zz_LsuPlugin_logic_flusher_cmdCounter;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_s0_remapped_1_exponent;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent;
  wire       [11:0]   _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_s0_remapped_4_exponent;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_s0_remapped_5_exponent;
  wire                _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_1;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_2;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_3;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_4;
  wire                _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_5;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_6;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_7;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_8;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_9;
  wire                _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_10;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_11;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_12;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_13;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_14;
  wire                _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_15;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_16;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_17;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_18;
  wire       [70:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_19;
  wire       [16:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_20;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_21;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_22;
  wire       [16:0]   _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_23;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_24;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_25;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent_1;
  wire       [53:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_1;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_2;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_3;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_4;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_5;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_6;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_7;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX;
  wire       [3:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_1;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_2;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_3;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_4;
  wire       [3:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_5;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_6;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_7;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_8;
  wire       [3:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_9;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_10;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_11;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_12;
  wire       [3:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_13;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_14;
  wire       [1:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_15;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_16;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_17;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_18;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_19;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_20;
  wire       [2:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_21;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_22;
  wire       [0:0]    _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_23;
  wire       [2:0]    _zz_65;
  reg        [2:0]    _zz_66;
  wire       [2:0]    _zz_67;
  reg        [2:0]    _zz_68;
  wire       [2:0]    _zz_69;
  wire       [1:0]    _zz_70;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_1;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_2;
  wire       [12:0]   _zz__zz_when_AFix_l1168_1_1;
  wire       [12:0]   _zz__zz_when_AFix_l1168_1_2;
  wire       [10:0]   _zz__zz_when_AFix_l1168_1_3;
  wire       [12:0]   _zz__zz_when_AFix_l1168_1_4;
  wire       [54:0]   _zz__zz_when_Utils_l1585_7;
  wire       [54:0]   _zz__zz_when_Utils_l1585_6;
  wire       [54:0]   _zz__zz_when_Utils_l1585_5;
  wire       [54:0]   _zz__zz_when_Utils_l1585_4;
  wire       [54:0]   _zz__zz_when_Utils_l1585_3;
  wire       [54:0]   _zz__zz_FpuPackerPlugin_logic_s1_subnormal_manShifter;
  wire       [54:0]   _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_2;
  wire       [54:0]   _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_3;
  wire       [0:0]    _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_4;
  wire       [1:0]    _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted;
  wire       [0:0]    _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted_1;
  wire       [29:0]   _zz_FpuPackerPlugin_logic_s1_incrBy;
  wire       [51:0]   _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry;
  wire       [52:0]   _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_1;
  wire       [30:0]   _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_2;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_2;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_3;
  wire       [1:0]    _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_4;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT_1;
  wire       [51:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_2;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_3;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_4;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_2;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_3;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_4;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX_1;
  wire       [11:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN;
  wire       [11:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_1;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_2;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_1;
  wire       [11:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_2;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_s2_fwb_value;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s0_VALUE_exponent;
  wire       [10:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL;
  wire       [12:0]   _zz_FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_3;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_2;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_3;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_1;
  wire       [31:0]   _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_2;
  wire       [9:0]    _zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK;
  wire       [15:0]   _zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK_1;
  wire       [3:0]    _zz__zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT_1;
  wire       [3:0]    _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed;
  wire       [1:0]    _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed_1;
  wire       [5:0]    _zz__zz_when_UInt_l128_1;
  wire       [2:0]    _zz__zz_when_UInt_l128_1_1;
  wire       [15:0]   _zz_PrefetcherRptPlugin_logic_storage_write_payload_data_address;
  wire       [4:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_1;
  wire       [4:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_2;
  wire       [4:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_3;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_2;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_3;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_4;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_5;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_6;
  wire       [11:0]   _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_7;
  wire       [4:0]    _zz_when_Prefetcher_l216;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_cached_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_io;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_3;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_2;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_3;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  wire                _zz_execute_lane0_api_hartsInflight;
  wire                _zz_execute_lane0_api_hartsInflight_1;
  wire                _zz_execute_lane0_api_hartsInflight_2;
  wire                _zz_execute_lane0_api_hartsInflight_3;
  wire       [0:0]    _zz_execute_lane0_api_hartsInflight_4;
  wire       [4:0]    _zz_execute_lane0_api_hartsInflight_5;
  wire                _zz_execute_lane0_api_hartsInflight_6;
  wire                _zz_execute_lane0_api_hartsInflight_7;
  wire                _zz_execute_lane0_api_hartsInflight_8;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS1_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_3;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_4;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_0_5;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS1_PHYS_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_0_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_0_3;
  wire                _zz_decode_ctrls_1_down_RS2_ENABLE_0_4;
  wire                _zz_decode_ctrls_1_down_RS2_ENABLE_0_5;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS2_PHYS_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_2;
  wire                _zz_decode_ctrls_1_down_RD_ENABLE_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0_4;
  wire       [10:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_8;
  wire                _zz_decode_ctrls_1_down_RD_ENABLE_0_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0_10;
  wire       [4:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_14;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_15;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_16;
  wire       [4:0]    _zz_decode_ctrls_1_down_RD_PHYS_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS3_ENABLE_0;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS3_PHYS_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_2;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_4;
  wire       [38:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_8;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_10;
  wire       [32:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_14;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_15;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_16;
  wire       [26:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_17;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_18;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_19;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_20;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_21;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_22;
  wire       [20:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_23;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_24;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_25;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_26;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_27;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_28;
  wire       [14:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_29;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_30;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_31;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_32;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_33;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_34;
  wire       [8:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_35;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_36;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_37;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_38;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_39;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_40;
  wire       [2:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_41;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire       [31:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS1_ENABLE_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_1_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_1_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_1_3;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_1_4;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS1_ENABLE_1_5;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS1_PHYS_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS2_ENABLE_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_1_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_1_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_1_3;
  wire                _zz_decode_ctrls_1_down_RS2_ENABLE_1_4;
  wire                _zz_decode_ctrls_1_down_RS2_ENABLE_1_5;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS2_PHYS_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_2;
  wire                _zz_decode_ctrls_1_down_RD_ENABLE_1_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_1_4;
  wire       [10:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_8;
  wire                _zz_decode_ctrls_1_down_RD_ENABLE_1_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_1_10;
  wire       [4:0]    _zz_decode_ctrls_1_down_RD_ENABLE_1_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_14;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_15;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_1_16;
  wire       [4:0]    _zz_decode_ctrls_1_down_RD_PHYS_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS3_ENABLE_1;
  wire       [4:0]    _zz_decode_ctrls_1_down_RS3_PHYS_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_2;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_4;
  wire       [38:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_8;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_10;
  wire       [32:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_14;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_15;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_16;
  wire       [26:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_17;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_18;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_19;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_20;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_21;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_22;
  wire       [20:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_23;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_24;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_25;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_26;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_27;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_28;
  wire       [14:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_29;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_30;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_31;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_32;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_33;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_34;
  wire       [8:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_35;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_36;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_37;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_1_38;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_1_39;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_40;
  wire       [2:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_1_41;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb;
  wire       [31:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5;
  reg        [0:0]    _zz_DispatchPlugin_logic_candidates_1_age;
  wire       [0:0]    _zz_DispatchPlugin_logic_candidates_1_age_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_candidates_2_age;
  wire       [1:0]    _zz_DispatchPlugin_logic_candidates_2_age_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_8;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_9;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_11;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_15;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_17;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_18;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_19;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_20;
  wire       [1:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_21;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_22;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_23;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_24;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_25;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_8;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_9;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_11;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_15;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_17;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_18;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_19;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_20;
  wire       [1:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_21;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_22;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_23;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_24;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_25;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_8;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_9;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_11;
  wire       [3:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_15;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_17;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_18;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_19;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_20;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_21;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_8;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_9;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_11;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_15;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_17;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_18;
  wire       [1:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_19;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_20;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_21;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_22;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_23;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_6;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_8;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_9;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_11;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_15;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_17;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_18;
  wire       [1:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_19;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_20;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_21;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_22;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_23;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_8;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_9;
  wire       [2:0]    _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_11;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_15;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_16;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_8;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_9;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_11;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_15;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_16;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_17;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_8;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_9;
  wire       [4:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_11;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_15;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_16;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_17;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_7;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_8;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_9;
  wire       [2:0]    _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_10;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_11;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_12;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_13;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_14;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_15;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_16;
  wire       [1:0]    _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [11:0]   _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [28:0]   _zz_BtbPlugin_logic_memWrite_payload_address;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent;
  wire       [51:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_1;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_2;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_1;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_2;
  wire       [11:0]   _zz_FpuUnpack_RS1_normalizer_exponent;
  wire       [11:0]   _zz_FpuUnpack_RS1_normalizer_exponent_1;
  wire       [6:0]    _zz_FpuUnpack_RS1_normalizer_exponent_2;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent;
  wire       [51:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_1;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_2;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_1;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_2;
  wire       [11:0]   _zz_FpuUnpack_RS2_normalizer_exponent;
  wire       [11:0]   _zz_FpuUnpack_RS2_normalizer_exponent_1;
  wire       [6:0]    _zz_FpuUnpack_RS2_normalizer_exponent_2;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent;
  wire       [51:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_1;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_2;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [10:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_1;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_2;
  wire       [11:0]   _zz_FpuUnpack_RS3_normalizer_exponent;
  wire       [11:0]   _zz_FpuUnpack_RS3_normalizer_exponent_1;
  wire       [6:0]    _zz_FpuUnpack_RS3_normalizer_exponent_2;
  wire       [31:0]   _zz_io_inputs_1_payload_data;
  wire       [5:0]    _zz_FpuUnpackerPlugin_logic_packPort_cmd_value_exponent;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_3;
  wire       [31:0]   _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3;
  wire       [3:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_2;
  wire       [4:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_16;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_17;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_18;
  wire       [4:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_19;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_3;
  wire       [31:0]   _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3;
  wire       [3:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_2;
  wire       [4:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_16;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_17;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_18;
  wire       [4:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_19;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0_1;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0_1;
  wire       [0:0]    _zz_FpuCmpPlugin_logic_iwb_payload;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_1;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_2;
  wire       [5:0]    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_3;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_4;
  wire       [53:0]   _zz__zz_when_Utils_l1585_2;
  wire       [53:0]   _zz__zz_when_Utils_l1585_1;
  wire       [53:0]   _zz__zz_when_Utils_l1585;
  wire       [53:0]   _zz__zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  wire       [53:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3;
  wire       [1:0]    _zz__zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6_1;
  wire       [53:0]   _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_2;
  wire       [31:0]   _zz_FpuF2iPlugin_logic_onResult_inverter;
  wire       [5:0]    _zz_FpuF2iPlugin_logic_onResult_expMax_1;
  wire       [5:0]    _zz_FpuF2iPlugin_logic_onResult_expMax_2;
  wire       [4:0]    _zz_FpuF2iPlugin_logic_onResult_expMax_3;
  wire       [5:0]    _zz_FpuF2iPlugin_logic_onResult_expMax_4;
  wire       [0:0]    _zz_FpuF2iPlugin_logic_onResult_expMax_5;
  wire       [5:0]    _zz_FpuF2iPlugin_logic_onResult_expMin;
  wire       [4:0]    _zz_FpuF2iPlugin_logic_onResult_expMin_1;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_overflow;
  wire       [6:0]    _zz_FpuF2iPlugin_logic_onResult_overflow_1;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_overflow_2;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_underflow;
  wire       [6:0]    _zz_FpuF2iPlugin_logic_onResult_underflow_1;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_underflow_2;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_underflow_3;
  wire       [11:0]   _zz_FpuF2iPlugin_logic_onResult_underflow_4;
  wire       [6:0]    _zz_FpuF2iPlugin_logic_onResult_underflow_5;
  wire       [11:0]   _zz_FpuAddPlugin_logic_addPort_cmd_rs1_exponent;
  wire       [11:0]   _zz_FpuAddPlugin_logic_addPort_cmd_rs2_exponent;
  wire       [12:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [12:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_1;
  wire       [12:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_2;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_3;
  wire       [12:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_4;
  wire       [11:0]   _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_5;
  wire       [110:0]  _zz_execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
  wire       [12:0]   _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0;
  wire       [12:0]   _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_1;
  wire       [12:0]   _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_2;
  wire       [12:0]   _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_3;
  wire       [1:0]    _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_4;
  wire       [104:0]  _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0;
  wire       [12:0]   _zz_FpuMulPlugin_logic_packPort_cmd_value_exponent;
  wire       [12:0]   _zz_FpuMulPlugin_logic_addPort_cmd_rs1_exponent;
  wire       [11:0]   _zz_FpuMulPlugin_logic_addPort_cmd_rs2_exponent;
  wire       [10:0]   _zz_FpuSqrtPlugin_logic_packPort_cmd_value_exponent;
  wire       [11:0]   _zz_FpuXxPlugin_logic_packPort_cmd_value_exponent;
  wire       [52:0]   _zz_early0_DivPlugin_logic_processing_a;
  wire       [52:0]   _zz_early0_DivPlugin_logic_processing_b;
  wire       [55:0]   _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0_1;
  wire       [53:0]   _zz_FpuDivPlugin_logic_onExecute_mantissa;
  wire       [0:0]    _zz_FpuDivPlugin_logic_onExecute_mantissa_1;
  wire       [12:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent;
  wire       [12:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent_1;
  wire       [12:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent_2;
  wire       [11:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent_3;
  wire       [12:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent_4;
  wire       [11:0]   _zz__zz_FpuDivPlugin_logic_onExecute_exponent_5;
  wire       [12:0]   _zz_FpuDivPlugin_logic_onExecute_exponent_1;
  wire       [12:0]   _zz_FpuDivPlugin_logic_onExecute_exponent_2;
  wire       [12:0]   _zz_FpuDivPlugin_logic_onExecute_exponent_3;
  wire       [1:0]    _zz_FpuDivPlugin_logic_onExecute_exponent_4;
  wire       [12:0]   _zz_FpuDivPlugin_logic_packPort_cmd_value_exponent;
  wire       [28:0]   _zz_BtbPlugin_logic_memWrite_payload_address_1;
  wire       [28:0]   _zz_BtbPlugin_logic_memRead_cmd_payload;
  wire       [30:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash;
  wire       [12:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_1;
  wire       [30:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_2;
  wire       [12:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_3;
  wire       [31:0]   _zz_BtbPlugin_logic_ras_write_payload_data;
  wire                _zz_AlignerPlugin_logic_buffer_flushIt;
  wire                _zz_AlignerPlugin_logic_buffer_flushIt_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_buffer_flushIt_2;
  wire       [1:0]    _zz_AlignerPlugin_logic_buffer_flushIt_3;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16;
  wire                _zz_DispatchPlugin_logic_candidates_0_cancel;
  wire                _zz_DispatchPlugin_logic_candidates_0_cancel_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_slotsFeeds_fit;
  wire       [1:0]    _zz_DispatchPlugin_logic_slotsFeeds_fit_1;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4;
  wire       [158:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2;
  wire       [152:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4;
  wire       [137:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5;
  wire       [15:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6;
  wire       [107:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8;
  wire       [70:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10;
  wire       [64:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11;
  wire       [7:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12;
  wire       [40:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15;
  wire       [158:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17;
  wire       [152:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19;
  wire       [137:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20;
  wire       [15:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21;
  wire       [107:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_22;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_23;
  wire       [70:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_24;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_25;
  wire       [64:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_26;
  wire       [7:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_27;
  wire       [40:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_28;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_29;
  wire       [0:0]    _zz_DispatchPlugin_logic_inserter_0_trap;
  wire       [0:0]    _zz_execute_ctrl0_up_LANE_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [3:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2;
  wire       [3:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_TRAP_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_RS3_ENABLE_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_DispatchPlugin_logic_inserter_1_trap;
  wire       [0:0]    _zz_execute_ctrl0_up_LANE_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2;
  wire       [1:0]    _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_TRAP_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_RS1_ENABLE_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_RS2_ENABLE_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_RD_ENABLE_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_RS3_ENABLE_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1;
  wire                _zz_decode_logic_flushes_0_onLanes_0_doIt;
  wire                _zz_decode_logic_flushes_0_onLanes_0_doIt_1;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_0_doIt_2;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_0_doIt_3;
  wire                _zz_decode_logic_flushes_0_onLanes_1_doIt;
  wire                _zz_decode_logic_flushes_0_onLanes_1_doIt_1;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_1_doIt_2;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_1_doIt_3;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_1;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_2;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_3;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_4;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_5;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_6;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt_7;
  wire       [3:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt_8;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_1;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_2;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_3;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt_4;
  wire       [2:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt_5;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [0:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1;
  wire       [31:0]   _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [2:0]    _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_self_pc;
  wire       [3:0]    _zz_PcPlugin_logic_harts_0_self_pc_1;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_6;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_7;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_8;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_9;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_10;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_11;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_12;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_13;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [2:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [1:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [1:0]    _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [2:0]    _zz_CsrRamPlugin_logic_flush_counter;
  wire       [0:0]    _zz_CsrRamPlugin_logic_flush_counter_1;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_1;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_3;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_4;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_5;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_6;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_7;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_8;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_9;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_10;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_11;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_12;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_13;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_14;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_15;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_1;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_3;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_4;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_5;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_6;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_7;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_8;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_9;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_10;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_11;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_12;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_13;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_14;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_15;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_1;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_2;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_3;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_4;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_5;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_6;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_7;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_8;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_9;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_10;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_11;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_12;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_13;
  wire                _zz_execute_ctrl1_down_float_RS1_lane0_14;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS1_lane0_15;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_1;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_2;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_3;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_4;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_5;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_6;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_7;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_8;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_9;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_10;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_11;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_12;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_13;
  wire                _zz_execute_ctrl1_down_float_RS2_lane0_14;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS2_lane0_15;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_1;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_2;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_3;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_4;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_5;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_6;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_7;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_8;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_9;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_10;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_11;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_12;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_13;
  wire                _zz_execute_ctrl1_down_float_RS3_lane0_14;
  wire       [63:0]   _zz_execute_ctrl1_down_float_RS3_lane0_15;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2;
  wire       [5:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_7;
  wire       [11:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_8;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_9;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_10;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_11;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_12;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_13;
  wire       [5:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_14;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_15;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_16;
  wire       [32:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_17;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_18;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_19;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_2;
  wire       [5:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_9;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_16;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_17;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_18;
  wire       [5:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_19;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1;
  wire       [32:0]   _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1;
  wire       [32:0]   _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2;
  wire                _zz_when_ExecuteLanePlugin_l306_2;
  wire                _zz_when_ExecuteLanePlugin_l306_2_1;
  wire                _zz_when_ExecuteLanePlugin_l306_2_2;
  wire                _zz_when_ExecuteLanePlugin_l306_2_3;
  wire       [0:0]    _zz_when_ExecuteLanePlugin_l306_2_4;
  wire       [0:0]    _zz_when_ExecuteLanePlugin_l306_2_5;
  wire                _zz_when_ExecuteLanePlugin_l306_4;
  wire                _zz_when_ExecuteLanePlugin_l306_4_1;
  wire       [31:0]   _zz_WhiteboxerPlugin_logic_csr_access_payload_address;
  wire                _zz_fetch_logic_flushes_0_doIt;
  wire                _zz_fetch_logic_flushes_0_doIt_1;
  wire       [0:0]    _zz_fetch_logic_flushes_0_doIt_2;
  wire       [1:0]    _zz_fetch_logic_flushes_0_doIt_3;
  wire                _zz_fetch_logic_flushes_1_doIt;
  wire                _zz_fetch_logic_flushes_1_doIt_1;
  wire       [0:0]    _zz_fetch_logic_flushes_1_doIt_2;
  wire       [0:0]    _zz_fetch_logic_flushes_1_doIt_3;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_1;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_3;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_4;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_5;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_6;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_7;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_8;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_9;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_10;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_11;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_12;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_13;
  wire                _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_14;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_15;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_1;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_3;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_4;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_5;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_6;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_7;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_8;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_9;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_10;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_11;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_12;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_13;
  wire                _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_14;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_15;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_2;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1;
  wire       [0:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2;
  wire                _zz_when_ExecuteLanePlugin_l306_7;
  wire                _zz_when_ExecuteLanePlugin_l306_7_1;
  wire                _zz_when_ExecuteLanePlugin_l306_7_2;
  wire                _zz_when_ExecuteLanePlugin_l306_7_3;
  wire                _zz_when_ExecuteLanePlugin_l306_7_4;
  wire                _zz_when_ExecuteLanePlugin_l306_7_5;
  wire                _zz_when_ExecuteLanePlugin_l306_7_6;
  wire                _zz_when_ExecuteLanePlugin_l306_9;
  wire                _zz_when_ExecuteLanePlugin_l306_9_1;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_loadExecute_data;
  wire                _zz_TrapPlugin_logic_initHold;
  wire                _zz_TrapPlugin_logic_initHold_1;
  wire                _zz_TrapPlugin_logic_initHold_2;
  reg        [1:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [2:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1;
  reg        [1:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  wire       [1:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1;
  wire       [11:0]   _zz_execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [11:0]   _zz_execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [11:0]   _zz_execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [11:0]   _zz_execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [11:0]   _zz_execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [11:0]   _zz_execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [11:0]   _zz_execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [12:0]   _zz_execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire                decode_ctrls_0_up_isValid;
  wire                fetch_logic_ctrls_0_up_isReady;
  wire                fetch_logic_ctrls_0_up_isValid;
  wire                execute_ctrl12_down_isReady;
  wire                execute_ctrl11_down_RD_ENABLE_lane0;
  reg        [63:0]   execute_ctrl12_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  reg        [0:0]    execute_ctrl12_up_LANE_AGE_lane0;
  reg        [4:0]    execute_ctrl12_up_RD_PHYS_lane0;
  reg        [0:0]    execute_ctrl12_up_RD_RFID_lane0;
  wire                execute_ctrl10_down_COMMIT_lane0;
  wire                execute_ctrl10_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl10_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl10_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl10_down_RD_ENABLE_lane0;
  wire       [15:0]   execute_ctrl10_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl10_down_TRAP_lane0;
  wire                execute_ctrl10_down_LANE_SEL_lane0;
  wire                execute_ctrl10_down_isReady;
  reg                 execute_ctrl11_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl11_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl11_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg        [0:0]    execute_ctrl11_up_LANE_AGE_lane0;
  reg        [4:0]    execute_ctrl11_up_RD_PHYS_lane0;
  reg        [0:0]    execute_ctrl11_up_RD_RFID_lane0;
  reg        [15:0]   execute_ctrl11_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl11_up_TRAP_lane0;
  wire                execute_ctrl9_down_COMMIT_lane0;
  wire                execute_ctrl9_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl9_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl9_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl9_down_RD_ENABLE_lane0;
  wire       [15:0]   execute_ctrl9_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl9_down_TRAP_lane0;
  wire                execute_ctrl9_down_LANE_SEL_lane0;
  wire                execute_ctrl9_down_isReady;
  reg        [63:0]   execute_ctrl10_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl10_up_COMMIT_lane0;
  reg                 execute_ctrl10_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl10_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl10_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl10_up_COMPLETED_lane0;
  reg        [0:0]    execute_ctrl10_up_LANE_AGE_lane0;
  reg        [4:0]    execute_ctrl10_up_RD_PHYS_lane0;
  reg        [0:0]    execute_ctrl10_up_RD_RFID_lane0;
  reg        [15:0]   execute_ctrl10_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl10_up_TRAP_lane0;
  wire                execute_ctrl8_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl8_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl8_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl8_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl8_down_RD_ENABLE_lane0;
  reg        [63:0]   execute_ctrl9_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl9_up_COMMIT_lane0;
  reg                 execute_ctrl9_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl9_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl9_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl9_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl9_up_COMPLETED_lane0;
  reg        [0:0]    execute_ctrl9_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl9_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl9_up_TRAP_lane0;
  wire                execute_ctrl7_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl7_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl7_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl7_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl7_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl7_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl7_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl7_down_RD_ENABLE_lane0;
  reg                 execute_ctrl8_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl8_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl8_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl8_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl8_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl8_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl8_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg        [0:0]    execute_ctrl8_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl8_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl8_up_TRAP_lane0;
  wire                execute_ctrl6_down_COMMIT_lane0;
  wire                execute_ctrl6_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl6_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl6_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl6_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl6_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl6_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl6_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl6_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl6_down_COMPLETION_AT_7_lane0;
  wire                execute_ctrl6_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl6_down_RD_ENABLE_lane0;
  wire       [15:0]   execute_ctrl6_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl6_down_TRAP_lane0;
  wire                execute_ctrl6_down_LANE_SEL_lane0;
  wire                execute_ctrl6_down_isReady;
  reg                 execute_ctrl7_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl7_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl7_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl7_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl7_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl7_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl7_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl7_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl7_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl7_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg        [0:0]    execute_ctrl7_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl7_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl7_up_TRAP_lane0;
  reg                 execute_ctrl7_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl5_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl5_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl5_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl5_down_BYPASSED_AT_7_lane0;
  wire                execute_ctrl5_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl5_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl5_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl5_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl5_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl5_down_COMPLETION_AT_7_lane0;
  wire                execute_ctrl5_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl5_down_RD_ENABLE_lane0;
  wire                execute_ctrl5_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  reg        [63:0]   execute_ctrl6_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl6_up_COMMIT_lane0;
  reg                 execute_ctrl6_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl6_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl6_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl6_up_BYPASSED_AT_7_lane0;
  reg                 execute_ctrl6_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl6_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl6_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl6_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl6_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl6_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl6_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl6_up_COMPLETED_lane0;
  reg        [0:0]    execute_ctrl6_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl6_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl6_up_TRAP_lane0;
  reg                 execute_ctrl6_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_logic_calc_SIGN_lane0;
  wire       [12:0]   execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [1:0]    execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode;
  wire                execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_quiet;
  wire                execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_sign;
  wire       [11:0]   execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mantissa;
  wire       [1:0]    execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode;
  wire                execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_quiet;
  wire                execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_sign;
  wire       [11:0]   execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mantissa;
  wire       [2:0]    execute_ctrl4_down_FpuUtils_ROUNDING_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_SUB2_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_SUB1_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_FMA_lane0;
  wire       [0:0]    execute_ctrl4_down_FpuUtils_FORMAT_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_7_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_6_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl4_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl4_down_COMPLETION_AT_5_lane0;
  wire                execute_ctrl4_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl4_down_COMPLETION_AT_7_lane0;
  wire                execute_ctrl4_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl4_down_FpuMulPlugin_SEL_lane0;
  reg        [105:0]  execute_ctrl5_up_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  reg        [12:0]   execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  reg        [31:0]   execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  reg        [31:0]   execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg        [1:0]    execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode;
  reg                 execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_quiet;
  reg                 execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_sign;
  reg        [11:0]   execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mantissa;
  reg        [1:0]    execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode;
  reg                 execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_quiet;
  reg                 execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_sign;
  reg        [11:0]   execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mantissa;
  reg        [1:0]    execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode;
  reg                 execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_quiet;
  reg                 execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_sign;
  reg        [11:0]   execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mantissa;
  reg        [2:0]    execute_ctrl5_up_FpuUtils_ROUNDING_lane0;
  reg                 execute_ctrl5_up_COMMIT_lane1;
  reg                 execute_ctrl5_up_FpuMulPlugin_SUB2_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_SUB1_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_FMA_lane0;
  reg        [0:0]    execute_ctrl5_up_FpuUtils_FORMAT_lane0;
  reg                 execute_ctrl5_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl5_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl5_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl5_up_BYPASSED_AT_7_lane0;
  reg                 execute_ctrl5_up_BYPASSED_AT_6_lane0;
  reg                 execute_ctrl5_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl5_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  reg                 execute_ctrl5_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl5_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl5_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl5_up_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl5_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl5_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl5_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl5_up_FpuMulPlugin_SEL_lane0;
  reg        [0:0]    execute_ctrl5_up_LANE_AGE_lane1;
  reg        [4:0]    execute_ctrl5_up_RD_PHYS_lane1;
  reg        [0:0]    execute_ctrl5_up_RD_RFID_lane1;
  reg        [0:0]    execute_ctrl5_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl5_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl5_up_TRAP_lane0;
  reg                 execute_ctrl5_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_logic_calc_SIGN_lane0;
  wire       [12:0]   execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [1:0]    execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode;
  wire                execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_quiet;
  wire                execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_sign;
  wire       [11:0]   execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mantissa;
  wire                execute_ctrl3_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  wire       [5:0]    execute_ctrl3_down_LsuPlugin_SB_PTR_lane0;
  wire       [11:0]   execute_ctrl3_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl3_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl3_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl3_down_LsuL1_CLEAN_lane0;
  wire       [7:0]    execute_ctrl3_down_LsuL1_MASK_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_WB_lane0;
  wire       [31:0]   execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire       [31:0]   execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire       [31:0]   execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire                execute_ctrl3_down_COMMIT_lane1;
  wire                execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  wire                execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  wire                execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  wire                execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  wire                execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  wire       [1:0]    execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [1:0]    execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1;
  wire                execute_ctrl3_down_SrcStageables_UNSIGNED_lane1;
  wire                execute_ctrl3_down_SrcStageables_ZERO_lane1;
  wire                execute_ctrl3_down_SrcStageables_REVERT_lane1;
  wire                execute_ctrl3_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                execute_ctrl3_down_COMPLETION_AT_4_lane1;
  wire                execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                execute_ctrl3_down_late1_BranchPlugin_SEL_lane1;
  wire                execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire                execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1;
  wire                execute_ctrl3_down_early1_BranchPlugin_SEL_lane1;
  wire       [1:0]    execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_SUB2_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_SUB1_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_FMA_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl3_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl3_down_MulPlugin_HIGH_lane0;
  wire       [1:0]    execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl3_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_7_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_6_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_5_lane0;
  wire       [1:0]    execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl3_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl3_down_SrcStageables_REVERT_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_5_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_7_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl3_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl3_down_FpuMulPlugin_SEL_lane0;
  wire                execute_ctrl3_down_FpuMvPlugin_SEL_FLOAT_lane0;
  wire                execute_ctrl3_down_FpuF2iPlugin_SEL_lane0;
  wire                execute_ctrl3_down_FpuCsrPlugin_DIRTY_lane0;
  wire                execute_ctrl3_down_late0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire                execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0;
  wire                execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl3_down_float_RS2_lane0;
  wire       [1:0]    execute_ctrl3_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl3_down_COMPLETED_lane1;
  wire       [15:0]   execute_ctrl3_down_Decode_UOP_ID_lane1;
  wire       [0:0]    execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [11:0]   execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [0:0]    execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0;
  reg                 execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  reg        [0:0]    execute_ctrl4_up_FpuF2iPlugin_logic_onShift_incrementPatched_lane0;
  reg                 execute_ctrl4_up_FpuF2iPlugin_logic_onShift_increment_lane0;
  reg                 execute_ctrl4_up_FpuF2iPlugin_logic_onShift_resign_lane0;
  reg        [53:0]   execute_ctrl4_up_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  reg                 execute_ctrl4_up_MMU_HAZARD_lane0;
  reg                 execute_ctrl4_up_MMU_REFILL_lane0;
  reg                 execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg        [31:0]   execute_ctrl4_up_MMU_TRANSLATED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  reg        [5:0]    execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  reg        [46:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [63:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [31:0]   execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [31:0]   execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  reg        [0:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  reg                 execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  reg        [12:0]   execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  reg        [1:0]    execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode;
  reg                 execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_quiet;
  reg                 execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_sign;
  reg        [11:0]   execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mantissa;
  reg        [1:0]    execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode;
  reg                 execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_quiet;
  reg                 execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_sign;
  reg        [11:0]   execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mantissa;
  reg        [1:0]    execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode;
  reg                 execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_quiet;
  reg                 execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_sign;
  reg        [11:0]   execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mantissa;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  reg        [63:0]   execute_ctrl4_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  reg        [5:0]    execute_ctrl4_up_LsuPlugin_SB_PTR_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl4_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl4_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl4_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl4_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl4_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1_SIZE_lane0;
  reg        [7:0]    execute_ctrl4_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_WB_lane0;
  reg        [2:0]    execute_ctrl4_up_FpuUtils_ROUNDING_lane0;
  reg        [31:0]   execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  reg        [31:0]   execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  reg        [31:0]   execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  reg        [31:0]   execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  reg        [31:0]   execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  reg        [31:0]   execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  reg        [5:0]    execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  reg        [22:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  reg        [22:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  reg        [39:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  reg        [39:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  reg        [56:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  reg        [56:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg        [7:0]    execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [63:0]   execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [31:0]   execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  reg                 execute_ctrl4_up_COMMIT_lane1;
  reg        [1:0]    execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 execute_ctrl4_up_SrcStageables_UNSIGNED_lane1;
  reg                 execute_ctrl4_up_SrcStageables_ZERO_lane1;
  reg                 execute_ctrl4_up_SrcStageables_REVERT_lane1;
  reg                 execute_ctrl4_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 execute_ctrl4_up_COMPLETION_AT_4_lane1;
  reg                 execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 execute_ctrl4_up_late1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1;
  reg                 execute_ctrl4_up_early1_BranchPlugin_SEL_lane1;
  reg        [1:0]    execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_SUB2_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_SUB1_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_FMA_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl4_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_LOAD_lane0;
  reg        [0:0]    execute_ctrl4_up_FpuUtils_FORMAT_lane0;
  reg                 execute_ctrl4_up_MulPlugin_HIGH_lane0;
  reg        [1:0]    execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 execute_ctrl4_up_SrcStageables_UNSIGNED_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_7_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_6_lane0;
  reg                 execute_ctrl4_up_BYPASSED_AT_5_lane0;
  reg        [1:0]    execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl4_up_SrcStageables_ZERO_lane0;
  reg                 execute_ctrl4_up_SrcStageables_REVERT_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_FpuMulPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_FpuMvPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl4_up_FpuF2iPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_FpuCsrPlugin_DIRTY_lane0;
  reg                 execute_ctrl4_up_late0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_early0_BranchPlugin_SEL_lane0;
  reg        [1:0]    execute_ctrl4_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    execute_ctrl4_up_LANE_AGE_lane1;
  reg        [4:0]    execute_ctrl4_up_RD_PHYS_lane1;
  reg        [0:0]    execute_ctrl4_up_RD_RFID_lane1;
  reg        [15:0]   execute_ctrl4_up_Decode_UOP_ID_lane1;
  reg                 execute_ctrl4_up_TRAP_lane1;
  reg        [31:0]   execute_ctrl4_up_PC_lane1;
  reg        [0:0]    execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   execute_ctrl4_up_Decode_UOP_lane1;
  reg        [0:0]    execute_ctrl4_up_LANE_AGE_lane0;
  reg        [15:0]   execute_ctrl4_up_Decode_UOP_ID_lane0;
  reg        [31:0]   execute_ctrl4_up_PC_lane0;
  reg                 execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  reg                 execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  reg        [0:0]    execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl4_up_Decode_UOP_lane0;
  wire                execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  wire                execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  wire                execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  wire                execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  wire                execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  wire       [1:0]    execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [0:0]    execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [1:0]    execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire                execute_ctrl2_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                execute_ctrl2_down_COMPLETION_AT_4_lane1;
  wire                execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                execute_ctrl2_down_late1_BranchPlugin_SEL_lane1;
  wire                execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire                execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1;
  wire       [1:0]    execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [0:0]    execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [1:0]    execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_SUB2_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_SUB1_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_FMA_lane0;
  wire                execute_ctrl2_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl2_down_MulPlugin_HIGH_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_7_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_6_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_5_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_4_lane0;
  wire       [1:0]    execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_8_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_5_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_3_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_11_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_7_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl2_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl2_down_FpuXxPlugin_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl2_down_FpuMvPlugin_SEL_INT_lane0;
  wire                execute_ctrl2_down_FpuMvPlugin_SEL_FLOAT_lane0;
  wire                execute_ctrl2_down_FpuF2iPlugin_SEL_lane0;
  wire                execute_ctrl2_down_FpuClassPlugin_SEL_lane0;
  wire                execute_ctrl2_down_FpuCsrPlugin_DIRTY_lane0;
  wire                execute_ctrl2_down_late0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire                execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0;
  wire                execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
  wire       [63:0]   execute_ctrl2_down_float_RS2_lane0;
  wire       [63:0]   execute_ctrl2_down_float_RS1_lane0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire                execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl2_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg                 execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  reg        [12:0]   execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  reg        [53:0]   execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  reg        [5:0]    execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  reg                 execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
  reg                 execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
  reg                 execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0;
  reg        [31:0]   execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  reg        [1:0]    execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode;
  reg                 execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_quiet;
  reg                 execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_sign;
  reg        [11:0]   execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mantissa;
  reg        [1:0]    execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode;
  reg                 execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_quiet;
  reg                 execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_sign;
  reg        [11:0]   execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mantissa;
  reg                 execute_ctrl3_up_FpuUnpack_RS1_badBoxing_HIT_lane0;
  reg        [1:0]    execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode;
  reg                 execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_quiet;
  reg                 execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_sign;
  reg        [11:0]   execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mantissa;
  reg                 execute_ctrl3_up_FpuUnpack_RS1_IS_SUBNORMAL_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  reg        [63:0]   execute_ctrl3_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  reg        [5:0]    execute_ctrl3_up_LsuPlugin_SB_PTR_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl3_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl3_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl3_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl3_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl3_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl3_up_LsuL1_SIZE_lane0;
  reg        [7:0]    execute_ctrl3_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_WB_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg        [2:0]    execute_ctrl3_up_FpuUtils_ROUNDING_lane0;
  reg        [31:0]   execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  reg        [31:0]   execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  reg        [31:0]   execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  reg        [31:0]   execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  reg        [5:0]    execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  reg        [22:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  reg        [22:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  reg        [39:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  reg        [39:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  reg        [56:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  reg        [56:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg        [7:0]    execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [63:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  reg                 execute_ctrl3_up_COMMIT_lane1;
  reg                 execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  reg                 execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  reg                 execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  reg                 execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  reg                 execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  reg                 execute_ctrl3_up_COMMIT_lane0;
  reg        [1:0]    execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  reg        [0:0]    execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  reg        [1:0]    execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 execute_ctrl3_up_SrcStageables_UNSIGNED_lane1;
  reg                 execute_ctrl3_up_SrcStageables_ZERO_lane1;
  reg                 execute_ctrl3_up_SrcStageables_REVERT_lane1;
  reg                 execute_ctrl3_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 execute_ctrl3_up_COMPLETION_AT_4_lane1;
  reg                 execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 execute_ctrl3_up_late1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1;
  reg                 execute_ctrl3_up_early1_BranchPlugin_SEL_lane1;
  reg        [1:0]    execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  reg        [0:0]    execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  reg        [1:0]    execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_SUB2_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_SUB1_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_FMA_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl3_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_LOAD_lane0;
  reg        [0:0]    execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0;
  reg        [0:0]    execute_ctrl3_up_FpuUtils_FORMAT_lane0;
  reg                 execute_ctrl3_up_MulPlugin_HIGH_lane0;
  reg        [1:0]    execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 execute_ctrl3_up_SrcStageables_UNSIGNED_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_7_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_6_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_5_lane0;
  reg                 execute_ctrl3_up_BYPASSED_AT_4_lane0;
  reg        [1:0]    execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl3_up_SrcStageables_ZERO_lane0;
  reg                 execute_ctrl3_up_SrcStageables_REVERT_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl3_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_FpuXxPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_FpuMulPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_FpuMvPlugin_SEL_INT_lane0;
  reg                 execute_ctrl3_up_FpuMvPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl3_up_FpuF2iPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_FpuCmpPlugin_SEL_CMP_lane0;
  reg                 execute_ctrl3_up_FpuCmpPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl3_up_FpuClassPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_FpuCsrPlugin_DIRTY_lane0;
  reg                 execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_late0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  reg        [1:0]    execute_ctrl3_up_AguPlugin_SIZE_lane0;
  reg                 execute_ctrl3_up_COMPLETED_lane1;
  reg        [0:0]    execute_ctrl3_up_LANE_AGE_lane1;
  reg        [4:0]    execute_ctrl3_up_RD_PHYS_lane1;
  reg        [0:0]    execute_ctrl3_up_RD_RFID_lane1;
  reg        [4:0]    execute_ctrl3_up_RS2_PHYS_lane1;
  reg        [0:0]    execute_ctrl3_up_RS2_RFID_lane1;
  reg        [4:0]    execute_ctrl3_up_RS1_PHYS_lane1;
  reg        [0:0]    execute_ctrl3_up_RS1_RFID_lane1;
  reg        [15:0]   execute_ctrl3_up_Decode_UOP_ID_lane1;
  reg                 execute_ctrl3_up_TRAP_lane1;
  reg        [31:0]   execute_ctrl3_up_PC_lane1;
  reg        [0:0]    execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   execute_ctrl3_up_Decode_UOP_lane1;
  reg        [0:0]    execute_ctrl3_up_LANE_AGE_lane0;
  reg        [4:0]    execute_ctrl3_up_RS2_PHYS_lane0;
  reg        [0:0]    execute_ctrl3_up_RS2_RFID_lane0;
  reg        [4:0]    execute_ctrl3_up_RS1_PHYS_lane0;
  reg        [0:0]    execute_ctrl3_up_RS1_RFID_lane0;
  reg        [15:0]   execute_ctrl3_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl3_up_TRAP_lane0;
  reg        [31:0]   execute_ctrl3_up_PC_lane0;
  reg                 execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  reg                 execute_ctrl3_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  reg        [0:0]    execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl3_up_Decode_UOP_lane0;
  wire       [1:0]    execute_ctrl1_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl1_down_COMPLETED_lane1;
  wire       [4:0]    execute_ctrl1_down_RD_PHYS_lane1;
  wire       [0:0]    execute_ctrl1_down_RD_RFID_lane1;
  wire       [15:0]   execute_ctrl1_down_Decode_UOP_ID_lane1;
  wire       [0:0]    execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [11:0]   execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1;
  wire                execute_ctrl1_down_COMPLETED_lane0;
  wire                execute_ctrl1_down_RS3_ENABLE_lane0;
  wire       [4:0]    execute_ctrl1_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl1_down_RD_RFID_lane0;
  wire                execute_ctrl1_down_RS2_ENABLE_lane0;
  wire                execute_ctrl1_down_RS1_ENABLE_lane0;
  wire       [15:0]   execute_ctrl1_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire       [0:0]    execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
  wire                execute_ctrl1_down_isReady;
  reg        [1:0]    execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  reg        [0:0]    execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  reg        [1:0]    execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 execute_ctrl2_up_SrcStageables_UNSIGNED_lane1;
  reg                 execute_ctrl2_up_BYPASSED_AT_3_lane1;
  reg                 execute_ctrl2_up_SrcStageables_ZERO_lane1;
  reg                 execute_ctrl2_up_SrcStageables_REVERT_lane1;
  reg        [1:0]    execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg                 execute_ctrl2_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 execute_ctrl2_up_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg                 execute_ctrl2_up_COMPLETION_AT_4_lane1;
  reg                 execute_ctrl2_up_COMPLETION_AT_2_lane1;
  reg                 execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_late1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_early1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1;
  reg        [1:0]    execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  reg        [0:0]    execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  reg        [1:0]    execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl2_up_FpuMulPlugin_SUB2_lane0;
  reg                 execute_ctrl2_up_FpuMulPlugin_SUB1_lane0;
  reg                 execute_ctrl2_up_FpuMulPlugin_FMA_lane0;
  reg                 execute_ctrl2_up_FpuAddPlugin_SUB_lane0;
  reg        [2:0]    execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl2_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_LOAD_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_EQUAL_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_LESS_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_SGNJ_RS1_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_INVERT_lane0;
  reg        [0:0]    execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0;
  reg        [0:0]    execute_ctrl2_up_FpuUtils_FORMAT_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  reg                 execute_ctrl2_up_DivPlugin_REM_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  reg                 execute_ctrl2_up_MulPlugin_HIGH_lane0;
  reg        [1:0]    execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_10_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_9_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_8_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_7_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_6_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_5_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_4_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_3_lane0;
  reg        [1:0]    execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl2_up_SrcStageables_ZERO_lane0;
  reg                 execute_ctrl2_up_SrcStageables_REVERT_lane0;
  reg        [1:0]    execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl2_up_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuUnpackerPlugin_SEL_I2F_lane0;
  reg                 execute_ctrl2_up_FpuDivPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuXxPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuSqrtPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuMulPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuAddPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuMvPlugin_SEL_INT_lane0;
  reg                 execute_ctrl2_up_FpuMvPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl2_up_FpuF2iPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_SEL_CMP_lane0;
  reg                 execute_ctrl2_up_FpuCmpPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl2_up_FpuClassPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_FpuCsrPlugin_DIRTY_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_late0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1;
  reg                 execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  reg        [31:0]   execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  reg        [1:0]    execute_ctrl2_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    execute_ctrl2_up_LANE_AGE_lane1;
  reg        [4:0]    execute_ctrl2_up_RS2_PHYS_lane1;
  reg        [0:0]    execute_ctrl2_up_RS2_RFID_lane1;
  reg        [4:0]    execute_ctrl2_up_RS1_PHYS_lane1;
  reg        [0:0]    execute_ctrl2_up_RS1_RFID_lane1;
  reg        [15:0]   execute_ctrl2_up_Decode_UOP_ID_lane1;
  reg        [31:0]   execute_ctrl2_up_PC_lane1;
  reg        [0:0]    execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   execute_ctrl2_up_Decode_UOP_lane1;
  reg        [0:0]    execute_ctrl2_up_LANE_AGE_lane0;
  reg        [0:0]    execute_ctrl2_up_RS3_RFID_lane0;
  reg        [4:0]    execute_ctrl2_up_RS2_PHYS_lane0;
  reg        [0:0]    execute_ctrl2_up_RS2_RFID_lane0;
  reg        [4:0]    execute_ctrl2_up_RS1_PHYS_lane0;
  reg        [0:0]    execute_ctrl2_up_RS1_RFID_lane0;
  reg        [15:0]   execute_ctrl2_up_Decode_UOP_ID_lane0;
  reg        [31:0]   execute_ctrl2_up_PC_lane0;
  reg                 execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  reg                 execute_ctrl2_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  reg        [0:0]    execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl2_up_Decode_UOP_lane0;
  wire       [0:0]    execute_ctrl0_down_lane1_LAYER_SEL_lane1;
  wire                execute_ctrl0_down_COMPLETED_lane1;
  wire       [4:0]    execute_ctrl0_down_RD_PHYS_lane1;
  wire       [0:0]    execute_ctrl0_down_RD_RFID_lane1;
  wire       [0:0]    execute_ctrl0_down_RS2_RFID_lane1;
  wire       [0:0]    execute_ctrl0_down_RS1_RFID_lane1;
  wire                execute_ctrl0_down_TRAP_lane1;
  wire       [31:0]   execute_ctrl0_down_PC_lane1;
  wire       [0:0]    execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [11:0]   execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   execute_ctrl0_down_Decode_UOP_lane1;
  wire       [0:0]    execute_ctrl0_down_lane0_LAYER_SEL_lane0;
  wire                execute_ctrl0_down_COMPLETED_lane0;
  wire       [0:0]    execute_ctrl0_down_RS3_RFID_lane0;
  wire                execute_ctrl0_down_RS3_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl0_down_RD_RFID_lane0;
  wire       [0:0]    execute_ctrl0_down_RS2_RFID_lane0;
  wire                execute_ctrl0_down_RS2_ENABLE_lane0;
  wire       [0:0]    execute_ctrl0_down_RS1_RFID_lane0;
  wire                execute_ctrl0_down_RS1_ENABLE_lane0;
  wire                execute_ctrl0_down_TRAP_lane0;
  wire       [31:0]   execute_ctrl0_down_PC_lane0;
  wire                execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  wire                execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl0_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire       [0:0]    execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
  reg        [1:0]    execute_ctrl1_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    execute_ctrl1_up_lane1_LAYER_SEL_lane1;
  reg                 execute_ctrl1_up_COMPLETED_lane1;
  reg        [0:0]    execute_ctrl1_up_LANE_AGE_lane1;
  reg        [4:0]    execute_ctrl1_up_RS2_PHYS_lane1;
  reg        [0:0]    execute_ctrl1_up_RS2_RFID_lane1;
  reg        [4:0]    execute_ctrl1_up_RS1_PHYS_lane1;
  reg        [0:0]    execute_ctrl1_up_RS1_RFID_lane1;
  reg        [15:0]   execute_ctrl1_up_Decode_UOP_ID_lane1;
  reg                 execute_ctrl1_up_TRAP_lane1;
  reg        [31:0]   execute_ctrl1_up_PC_lane1;
  reg        [0:0]    execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   execute_ctrl1_up_Decode_UOP_lane1;
  reg        [0:0]    execute_ctrl1_up_lane0_LAYER_SEL_lane0;
  reg                 execute_ctrl1_up_COMPLETED_lane0;
  reg        [0:0]    execute_ctrl1_up_LANE_AGE_lane0;
  reg        [4:0]    execute_ctrl1_up_RS3_PHYS_lane0;
  reg        [0:0]    execute_ctrl1_up_RS3_RFID_lane0;
  reg                 execute_ctrl1_up_RS3_ENABLE_lane0;
  reg        [4:0]    execute_ctrl1_up_RS2_PHYS_lane0;
  reg        [0:0]    execute_ctrl1_up_RS2_RFID_lane0;
  reg                 execute_ctrl1_up_RS2_ENABLE_lane0;
  reg        [4:0]    execute_ctrl1_up_RS1_PHYS_lane0;
  reg        [0:0]    execute_ctrl1_up_RS1_RFID_lane0;
  reg                 execute_ctrl1_up_RS1_ENABLE_lane0;
  reg        [15:0]   execute_ctrl1_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl1_up_TRAP_lane0;
  reg        [31:0]   execute_ctrl1_up_PC_lane0;
  reg                 execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  reg                 execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  reg                 execute_ctrl1_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  reg                 execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  reg        [0:0]    execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl1_up_Decode_UOP_lane0;
  wire                decode_ctrls_1_down_isReady;
  wire                decode_ctrls_0_down_Prediction_ALIGN_REDO_1;
  wire       [3:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [3:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [31:0]   decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1;
  wire                decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1;
  wire       [11:0]   decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [0:0]    decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1;
  wire                decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_1;
  wire                decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
  wire       [3:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [3:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
  wire       [11:0]   decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [0:0]    decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_down_isValid;
  wire                decode_ctrls_0_down_isReady;
  reg                 decode_ctrls_1_up_Prediction_ALIGN_REDO_1;
  reg        [3:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  reg        [3:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  reg        [31:0]   decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1;
  reg                 decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1;
  reg        [11:0]   decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3;
  reg        [9:0]    decode_ctrls_1_up_Decode_DOP_ID_1;
  reg        [31:0]   decode_ctrls_1_up_PC_1;
  reg        [0:0]    decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1;
  reg                 decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_1;
  reg                 decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  reg        [3:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  reg        [3:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  reg        [31:0]   decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  reg                 decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  reg        [11:0]   decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3;
  reg        [9:0]    decode_ctrls_1_up_Decode_DOP_ID_0;
  reg        [31:0]   decode_ctrls_1_up_PC_0;
  reg        [0:0]    decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  reg                 decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_0;
  wire       [9:0]    fetch_logic_ctrls_1_down_Fetch_ID;
  wire                fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_1_down_isValid;
  wire                fetch_logic_ctrls_1_down_isReady;
  reg                 fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  reg                 fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  reg                 fetch_logic_ctrls_2_up_MMU_HAZARD;
  reg                 fetch_logic_ctrls_2_up_MMU_REFILL;
  reg        [3:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  reg        [3:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  reg        [31:0]   fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  reg        [1:0]    fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE;
  reg                 fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  reg        [31:0]   fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  reg        [63:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  reg        [63:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  reg        [0:0]    fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg        [11:0]   fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  reg        [9:0]    fetch_logic_ctrls_2_up_Fetch_ID;
  reg                 fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_0_down_isValid;
  reg        [1:0]    fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  reg                 fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3;
  reg        [11:0]   fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  reg        [5:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  reg        [0:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg        [9:0]    fetch_logic_ctrls_1_up_Fetch_ID;
  reg                 fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_2_up_valid;
  wire                decode_ctrls_1_down_valid;
  reg                 fetch_logic_ctrls_1_down_valid;
  wire                decode_ctrls_0_down_valid;
  reg                 fetch_logic_ctrls_0_down_valid;
  wire                execute_ctrl0_up_ready;
  wire                execute_ctrl0_down_ready;
  wire                execute_ctrl1_up_ready;
  wire                execute_ctrl1_down_ready;
  wire                execute_ctrl2_up_ready;
  wire                execute_ctrl2_down_ready;
  wire                execute_ctrl3_up_ready;
  wire                execute_ctrl3_down_ready;
  wire                execute_ctrl4_up_ready;
  wire                execute_ctrl4_down_ready;
  wire                execute_ctrl5_up_ready;
  wire                execute_ctrl5_down_ready;
  wire                execute_ctrl6_up_ready;
  wire                execute_ctrl6_down_ready;
  wire                execute_ctrl7_up_ready;
  wire                execute_ctrl7_down_ready;
  wire                execute_ctrl8_up_ready;
  wire                execute_ctrl8_down_ready;
  wire                execute_ctrl9_up_ready;
  wire                execute_ctrl9_down_ready;
  wire                execute_ctrl10_up_ready;
  wire                execute_ctrl10_down_ready;
  wire                fetch_logic_ctrls_0_down_ready;
  wire                execute_ctrl11_up_ready;
  wire                decode_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_1_up_cancel;
  wire                execute_ctrl11_down_ready;
  reg                 decode_ctrls_0_down_ready;
  wire                fetch_logic_ctrls_1_down_ready;
  wire                execute_ctrl12_up_ready;
  wire                fetch_logic_ctrls_2_up_ready;
  wire                fetch_logic_ctrls_2_up_cancel;
  wire                execute_ctrl4_down_AguPlugin_ATOMIC_lane0;
  wire       [31:0]   execute_ctrl4_down_MMU_TRANSLATED_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl4_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl12_down_ready;
  reg                 execute_ctrl2_up_TRAP_lane1;
  wire                execute_ctrl2_up_COMMIT_lane1;
  wire                execute_ctrl3_down_TRAP_lane1;
  wire       [0:0]    execute_ctrl5_down_LANE_AGE_lane1;
  wire                execute_ctrl4_down_RD_ENABLE_lane1;
  reg                 execute_ctrl4_RD_ENABLE_lane1_bypass;
  reg                 execute_ctrl4_LANE_SEL_lane1_bypass;
  wire                execute_ctrl3_down_RD_ENABLE_lane1;
  reg                 execute_ctrl3_RD_ENABLE_lane1_bypass;
  wire                execute_ctrl3_down_LANE_SEL_lane1;
  reg                 execute_ctrl3_LANE_SEL_lane1_bypass;
  wire       [0:0]    execute_ctrl3_down_LANE_AGE_lane1;
  wire                execute_ctrl2_down_RD_ENABLE_lane1;
  reg                 execute_ctrl2_RD_ENABLE_lane1_bypass;
  reg                 execute_ctrl2_LANE_SEL_lane1_bypass;
  wire                execute_ctrl1_down_RD_ENABLE_lane1;
  reg                 execute_ctrl1_RD_ENABLE_lane1_bypass;
  wire                execute_ctrl1_down_LANE_SEL_lane1;
  reg                 execute_ctrl1_LANE_SEL_lane1_bypass;
  wire       [0:0]    execute_ctrl1_down_LANE_AGE_lane1;
  wire                execute_ctrl0_down_RD_ENABLE_lane1;
  reg                 execute_ctrl0_RD_ENABLE_lane1_bypass;
  reg                 execute_ctrl0_LANE_SEL_lane1_bypass;
  wire       [0:0]    execute_ctrl0_down_LANE_AGE_lane1;
  wire                execute_ctrl1_down_TRAP_lane1;
  wire       [1:0]    execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [0:0]    execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [1:0]    execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [1:0]    execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
  wire                execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
  wire                execute_ctrl1_down_BYPASSED_AT_3_lane1;
  wire                execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1;
  wire                execute_ctrl1_down_SrcStageables_ZERO_lane1;
  wire                execute_ctrl1_down_SrcStageables_REVERT_lane1;
  wire       [1:0]    execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg                 execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg                 execute_ctrl1_down_COMPLETION_AT_4_lane1;
  reg                 execute_ctrl1_down_COMPLETION_AT_2_lane1;
  reg                 execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
  reg                 execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    execute_ctrl1_down_lane1_LAYER_SEL_lane1;
  wire                execute_ctrl4_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                execute_ctrl2_down_TRAP_lane1;
  wire                execute_ctrl2_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg        [31:0]   execute_ctrl3_up_integer_RS2_lane1;
  wire       [31:0]   execute_ctrl3_integer_RS2_lane1_bypass;
  wire       [0:0]    execute_ctrl3_down_RS2_RFID_lane1;
  wire       [4:0]    execute_ctrl3_down_RS2_PHYS_lane1;
  reg        [31:0]   execute_ctrl2_up_integer_RS2_lane1;
  wire       [31:0]   execute_ctrl2_down_integer_RS2_lane1;
  wire       [31:0]   execute_ctrl2_integer_RS2_lane1_bypass;
  wire       [0:0]    execute_ctrl2_down_RS2_RFID_lane1;
  wire       [4:0]    execute_ctrl2_down_RS2_PHYS_lane1;
  wire       [0:0]    execute_ctrl1_down_RS2_RFID_lane1;
  wire       [4:0]    execute_ctrl1_down_RS2_PHYS_lane1;
  wire       [4:0]    execute_ctrl0_down_RS2_PHYS_lane1;
  reg        [31:0]   execute_ctrl3_up_integer_RS1_lane1;
  wire       [31:0]   execute_ctrl3_integer_RS1_lane1_bypass;
  wire       [0:0]    execute_ctrl3_down_RS1_RFID_lane1;
  wire       [4:0]    execute_ctrl3_down_RS1_PHYS_lane1;
  reg        [31:0]   execute_ctrl2_up_integer_RS1_lane1;
  wire       [31:0]   execute_ctrl2_down_integer_RS1_lane1;
  wire       [31:0]   execute_ctrl2_integer_RS1_lane1_bypass;
  wire       [0:0]    execute_ctrl2_down_RS1_RFID_lane1;
  wire       [4:0]    execute_ctrl2_down_RS1_PHYS_lane1;
  wire       [0:0]    execute_ctrl1_down_RS1_RFID_lane1;
  wire       [4:0]    execute_ctrl1_down_RS1_PHYS_lane1;
  wire       [0:0]    execute_ctrl12_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl11_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl10_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl9_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl8_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl7_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl6_down_LANE_AGE_lane0;
  wire       [0:0]    execute_ctrl5_down_LANE_AGE_lane0;
  wire                execute_ctrl4_down_RD_ENABLE_lane0;
  reg                 execute_ctrl4_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl4_LANE_SEL_lane0_bypass;
  wire                execute_ctrl3_down_RD_ENABLE_lane0;
  reg                 execute_ctrl3_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl3_LANE_SEL_lane0_bypass;
  wire       [0:0]    execute_ctrl3_down_LANE_AGE_lane0;
  wire                execute_ctrl2_down_RD_ENABLE_lane0;
  reg                 execute_ctrl2_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl2_LANE_SEL_lane0_bypass;
  wire                execute_ctrl1_down_RD_ENABLE_lane0;
  reg                 execute_ctrl1_RD_ENABLE_lane0_bypass;
  wire                execute_ctrl1_down_LANE_SEL_lane0;
  reg                 execute_ctrl1_LANE_SEL_lane0_bypass;
  wire       [0:0]    execute_ctrl1_down_LANE_AGE_lane0;
  wire                execute_ctrl0_down_RD_ENABLE_lane0;
  reg                 execute_ctrl0_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl0_LANE_SEL_lane0_bypass;
  wire       [0:0]    execute_ctrl0_down_LANE_AGE_lane0;
  wire                execute_ctrl1_down_TRAP_lane0;
  wire       [1:0]    execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [0:0]    execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [1:0]    execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0;
  wire                execute_ctrl1_down_FpuMulPlugin_SUB2_lane0;
  wire                execute_ctrl1_down_FpuMulPlugin_SUB1_lane0;
  wire                execute_ctrl1_down_FpuMulPlugin_FMA_lane0;
  wire                execute_ctrl1_down_FpuAddPlugin_SUB_lane0;
  wire       [2:0]    execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire                execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire                execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire                execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0;
  wire                execute_ctrl1_down_FpuCmpPlugin_LESS_lane0;
  wire                execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0;
  wire                execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0;
  wire       [0:0]    execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0;
  wire       [0:0]    execute_ctrl1_down_FpuUtils_FORMAT_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl1_down_DivPlugin_REM_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire                execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [1:0]    execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_10_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_9_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_8_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_7_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_6_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_5_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_4_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire       [1:0]    execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0;
  reg                 execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0;
  reg                 execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0;
  reg                 execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0;
  reg                 execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0;
  reg                 execute_ctrl1_down_FpuDivPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuXxPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuMulPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuAddPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl1_down_AguPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0;
  reg                 execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl1_down_FpuF2iPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0;
  reg                 execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0;
  reg                 execute_ctrl1_down_FpuClassPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0;
  reg                 execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    execute_ctrl1_down_lane0_LAYER_SEL_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
  wire                execute_ctrl8_down_TRAP_lane0;
  wire                execute_ctrl8_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                execute_ctrl5_down_TRAP_lane0;
  wire                execute_ctrl5_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  wire                execute_ctrl3_down_TRAP_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  wire                execute_ctrl11_down_TRAP_lane0;
  wire                execute_ctrl11_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl7_down_TRAP_lane0;
  wire                execute_ctrl7_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire       [63:0]   execute_ctrl1_down_float_RS3_lane0;
  wire       [0:0]    execute_ctrl1_down_RS3_RFID_lane0;
  wire       [4:0]    execute_ctrl1_down_RS3_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS3_PHYS_lane0;
  wire       [63:0]   execute_ctrl1_down_float_RS2_lane0;
  wire       [63:0]   execute_ctrl1_down_float_RS1_lane0;
  wire       [63:0]   execute_ctrl12_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [0:0]    execute_ctrl12_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl12_down_RD_PHYS_lane0;
  reg                 execute_ctrl12_up_RD_ENABLE_lane0;
  reg                 execute_ctrl12_up_LANE_SEL_lane0;
  wire       [0:0]    execute_ctrl11_down_RD_RFID_lane0;
  wire       [0:0]    execute_ctrl10_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl10_down_RD_PHYS_lane0;
  reg                 execute_ctrl10_up_RD_ENABLE_lane0;
  wire       [0:0]    execute_ctrl9_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl9_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl8_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl8_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl7_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl7_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl6_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl6_down_RD_PHYS_lane0;
  reg        [31:0]   execute_ctrl3_up_integer_RS2_lane0;
  wire       [31:0]   execute_ctrl3_integer_RS2_lane0_bypass;
  wire       [0:0]    execute_ctrl3_down_RS2_RFID_lane0;
  wire       [4:0]    execute_ctrl3_down_RS2_PHYS_lane0;
  wire       [31:0]   execute_ctrl2_down_integer_RS2_lane0;
  wire       [31:0]   execute_ctrl2_integer_RS2_lane0_bypass;
  wire       [4:0]    execute_ctrl2_down_RS2_PHYS_lane0;
  wire       [0:0]    execute_ctrl1_down_RS2_RFID_lane0;
  wire       [4:0]    execute_ctrl1_down_RS2_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS2_PHYS_lane0;
  reg        [31:0]   execute_ctrl3_up_integer_RS1_lane0;
  wire       [31:0]   execute_ctrl3_integer_RS1_lane0_bypass;
  wire       [0:0]    execute_ctrl3_down_RS1_RFID_lane0;
  wire       [4:0]    execute_ctrl3_down_RS1_PHYS_lane0;
  wire       [31:0]   execute_ctrl2_down_integer_RS1_lane0;
  wire       [31:0]   execute_ctrl2_integer_RS1_lane0_bypass;
  wire       [4:0]    execute_ctrl2_down_RS1_PHYS_lane0;
  wire       [31:0]   execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [0:0]    execute_ctrl5_down_RD_RFID_lane1;
  wire       [4:0]    execute_ctrl5_down_RD_PHYS_lane1;
  reg                 execute_ctrl5_up_RD_ENABLE_lane1;
  reg                 execute_ctrl5_up_LANE_SEL_lane1;
  wire       [0:0]    execute_ctrl5_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl5_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl4_down_RD_RFID_lane1;
  wire       [0:0]    execute_ctrl4_down_RD_RFID_lane0;
  wire       [0:0]    execute_ctrl3_down_RD_RFID_lane1;
  wire       [4:0]    execute_ctrl3_down_RD_PHYS_lane1;
  reg                 execute_ctrl3_up_RD_ENABLE_lane1;
  wire       [0:0]    execute_ctrl3_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl3_down_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl2_down_RD_RFID_lane1;
  wire       [4:0]    execute_ctrl2_down_RD_PHYS_lane1;
  wire       [0:0]    execute_ctrl1_down_RS1_RFID_lane0;
  wire       [0:0]    execute_ctrl2_down_RD_RFID_lane0;
  wire       [4:0]    execute_ctrl1_down_RS1_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS1_PHYS_lane0;
  reg                 _zz_1;
  wire                execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
  wire                execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0;
  wire                fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
  wire                fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
  wire                fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE;
  wire                fetch_logic_ctrls_1_down_MMU_ALLOW_READ;
  wire                fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
  wire                fetch_logic_ctrls_1_down_MMU_HAZARD;
  wire                fetch_logic_ctrls_1_down_MMU_REFILL;
  wire                execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  wire       [4:0]    execute_ctrl2_down_RD_PHYS_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
  wire                fetch_logic_ctrls_0_up_isFiring;
  reg        [9:0]    fetch_logic_ctrls_0_up_Fetch_ID;
  wire                fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  wire       [31:0]   fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_0_up_valid;
  reg                 PcPlugin_logic_harts_0_aggregator_fault_1;
  reg        [31:0]   PcPlugin_logic_harts_0_aggregator_target_1;
  wire       [0:0]    execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [0:0]    execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire                execute_ctrl4_down_TRAP_lane1;
  wire                execute_ctrl5_down_COMMIT_lane1;
  wire                execute_ctrl5_down_LANE_SEL_lane1;
  wire       [4:0]    execute_ctrl0_down_RS1_PHYS_lane1;
  wire                decode_ctrls_0_down_TRAP_1;
  wire                decode_ctrls_0_down_TRAP_0;
  wire                decode_ctrls_1_down_LANE_SEL_1;
  reg                 decode_ctrls_1_LANE_SEL_1_bypass;
  wire                decode_ctrls_1_down_LANE_SEL_0;
  reg                 decode_ctrls_1_LANE_SEL_0_bypass;
  wire                decode_ctrls_0_down_LANE_SEL_1;
  reg                 decode_ctrls_0_LANE_SEL_1_bypass;
  wire                decode_ctrls_0_down_LANE_SEL_0;
  reg                 decode_ctrls_0_LANE_SEL_0_bypass;
  wire       [0:0]    execute_ctrl0_up_lane1_LAYER_SEL_lane1;
  wire                execute_ctrl0_up_COMPLETED_lane1;
  wire       [0:0]    execute_ctrl0_up_LANE_AGE_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1;
  wire       [4:0]    execute_ctrl0_up_RS3_PHYS_lane1;
  wire       [0:0]    execute_ctrl0_up_RS3_RFID_lane1;
  wire                execute_ctrl0_up_RS3_ENABLE_lane1;
  wire       [4:0]    execute_ctrl0_up_RD_PHYS_lane1;
  wire       [0:0]    execute_ctrl0_up_RD_RFID_lane1;
  reg                 execute_ctrl0_up_RD_ENABLE_lane1;
  wire       [4:0]    execute_ctrl0_up_RS2_PHYS_lane1;
  wire       [0:0]    execute_ctrl0_up_RS2_RFID_lane1;
  wire                execute_ctrl0_up_RS2_ENABLE_lane1;
  wire       [4:0]    execute_ctrl0_up_RS1_PHYS_lane1;
  wire       [0:0]    execute_ctrl0_up_RS1_RFID_lane1;
  wire                execute_ctrl0_up_RS1_ENABLE_lane1;
  wire       [15:0]   execute_ctrl0_up_Decode_UOP_ID_lane1;
  wire                execute_ctrl0_up_TRAP_lane1;
  wire       [31:0]   execute_ctrl0_up_PC_lane1;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane1;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane1;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane1;
  wire                execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane1;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane1;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane1;
  wire                execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane1;
  wire       [0:0]    execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1;
  reg                 execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1;
  wire                execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1;
  wire       [11:0]   execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   execute_ctrl0_up_Decode_UOP_lane1;
  wire                execute_ctrl0_up_LANE_SEL_lane1;
  wire       [0:0]    execute_ctrl0_up_lane0_LAYER_SEL_lane0;
  wire                execute_ctrl0_up_COMPLETED_lane0;
  wire       [0:0]    execute_ctrl0_up_LANE_AGE_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [4:0]    execute_ctrl0_up_RS3_PHYS_lane0;
  wire       [0:0]    execute_ctrl0_up_RS3_RFID_lane0;
  wire                execute_ctrl0_up_RS3_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RD_PHYS_lane0;
  wire       [0:0]    execute_ctrl0_up_RD_RFID_lane0;
  reg                 execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS2_PHYS_lane0;
  wire       [0:0]    execute_ctrl0_up_RS2_RFID_lane0;
  wire                execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS1_PHYS_lane0;
  wire       [0:0]    execute_ctrl0_up_RS1_RFID_lane0;
  wire                execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [15:0]   execute_ctrl0_up_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_up_TRAP_lane0;
  wire       [31:0]   execute_ctrl0_up_PC_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane0;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire                execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane0;
  wire       [0:0]    execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  reg                 execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [11:0]   execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl0_up_Decode_UOP_lane0;
  wire                execute_ctrl0_up_LANE_SEL_lane0;
  wire                decode_ctrls_0_up_isMoving;
  reg        [3:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
  reg        [3:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  wire       [31:0]   fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
  wire       [1:0]    fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE;
  wire                fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
  wire                fetch_logic_ctrls_1_up_isCancel;
  wire                fetch_logic_ctrls_1_up_isReady;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
  (* keep , syn_keep *) wire       [11:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [30:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  wire       [1:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire                fetch_logic_ctrls_1_up_isValid;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  (* keep , syn_keep *) wire       [11:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [30:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire       [15:0]   execute_ctrl0_down_Decode_UOP_ID_lane1;
  wire                execute_ctrl0_down_LANE_SEL_lane1;
  wire       [15:0]   execute_ctrl0_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_down_isReady;
  wire                execute_ctrl0_down_LANE_SEL_lane0;
  wire       [9:0]    decode_ctrls_1_down_Decode_DOP_ID_1;
  wire       [9:0]    decode_ctrls_1_down_Decode_DOP_ID_0;
  wire       [55:0]   execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0;
  wire                execute_ctrl2_down_FpuDivPlugin_SEL_lane0;
  wire                execute_ctrl3_down_FpuXxPlugin_SEL_lane0;
  wire                execute_ctrl2_down_FpuSqrtPlugin_SEL_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_SUB2_lane0;
  wire       [1:0]    execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode;
  wire                execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_quiet;
  wire                execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_sign;
  wire       [11:0]   execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mantissa;
  wire                execute_ctrl5_down_FpuMulPlugin_SUB1_lane0;
  wire       [2:0]    execute_ctrl5_down_FpuUtils_ROUNDING_lane0;
  wire       [0:0]    execute_ctrl5_down_FpuUtils_FORMAT_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_logic_calc_SIGN_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_FMA_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_SEL_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  wire       [1:0]    execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode;
  wire                execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_quiet;
  wire                execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_sign;
  wire       [11:0]   execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mantissa;
  wire       [1:0]    execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode;
  wire                execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_quiet;
  wire                execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_sign;
  wire       [11:0]   execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mantissa;
  wire                execute_ctrl5_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  wire                execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  wire       [104:0]  execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0;
  wire       [12:0]   execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0;
  wire       [12:0]   execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire       [105:0]  execute_ctrl5_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
  wire       [105:0]  execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_SEL_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  wire                execute_ctrl2_down_FpuMulPlugin_logic_calc_SIGN_lane0;
  wire       [12:0]   execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  wire                execute_ctrl2_down_FpuAddPlugin_SUB_lane0;
  wire                execute_ctrl2_down_FpuAddPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_FpuF2iPlugin_logic_onResult_RESULT_lane0;
  reg                 execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NX_lane0;
  reg                 execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NV_lane0;
  wire                execute_ctrl4_down_FpuF2iPlugin_logic_onShift_increment_lane0;
  wire       [1:0]    execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode;
  wire                execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_quiet;
  wire                execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign;
  wire       [11:0]   execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mantissa;
  wire       [0:0]    execute_ctrl4_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0;
  wire                execute_ctrl4_down_FpuF2iPlugin_logic_onShift_resign_lane0;
  wire                execute_ctrl4_down_FpuF2iPlugin_SEL_lane0;
  wire       [53:0]   execute_ctrl4_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  wire       [0:0]    execute_ctrl3_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0;
  wire                execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0;
  wire       [2:0]    execute_ctrl3_down_FpuUtils_ROUNDING_lane0;
  wire                execute_ctrl3_down_FpuF2iPlugin_logic_onShift_resign_lane0;
  wire       [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2;
  reg        [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1;
  wire       [5:0]    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  wire       [53:0]   execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  wire       [53:0]   execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  reg        [53:0]   _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  reg        [53:0]   _zz_when_Utils_l1585;
  reg        [53:0]   _zz_when_Utils_l1585_1;
  reg        [53:0]   _zz_when_Utils_l1585_2;
  wire       [5:0]    execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  wire       [11:0]   execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0;
  wire                execute_ctrl3_down_FpuUnpack_RS1_badBoxing_HIT_lane0;
  wire                execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
  wire       [1:0]    execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode;
  wire                execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_quiet;
  wire                execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_sign;
  wire       [11:0]   execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mantissa;
  reg        [63:0]   execute_ctrl3_up_float_RS2_lane0;
  wire                execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0;
  wire       [0:0]    execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0;
  wire                execute_ctrl3_down_FpuCmpPlugin_SEL_FLOAT_lane0;
  wire                execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
  wire                execute_ctrl3_down_FpuCmpPlugin_SEL_CMP_lane0;
  wire       [0:0]    execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_SEL_FLOAT_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_INVERT_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_SGNJ_RS1_lane0;
  reg                 execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_EQUAL_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1MantissaSmaller_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0;
  reg                 execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1Equal_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_bothZero_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_NV_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_LESS_lane0;
  wire                execute_ctrl2_down_FpuCmpPlugin_SEL_CMP_lane0;
  wire                execute_ctrl3_down_FpuClassPlugin_SEL_lane0;
  wire                execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0;
  wire       [1:0]    execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode;
  wire                execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet;
  wire                execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign;
  wire       [11:0]   execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent;
  wire       [51:0]   execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mantissa;
  wire       [0:0]    execute_ctrl3_down_FpuUtils_FORMAT_lane0;
  wire       [4:0]    execute_ctrl11_down_RD_PHYS_lane0;
  wire                execute_ctrl11_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire       [15:0]   execute_ctrl11_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl11_down_COMMIT_lane0;
  reg                 execute_ctrl11_up_RD_ENABLE_lane0;
  wire                execute_ctrl11_down_isReady;
  wire                execute_ctrl11_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl11_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl11_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [15:0]   execute_ctrl8_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl8_down_COMMIT_lane0;
  wire                execute_ctrl8_down_isReady;
  wire                execute_ctrl8_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl8_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl8_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [15:0]   execute_ctrl7_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl7_down_COMMIT_lane0;
  wire                execute_ctrl7_down_isReady;
  wire                execute_ctrl7_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl7_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl7_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [15:0]   execute_ctrl5_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl5_down_COMMIT_lane0;
  wire                execute_ctrl5_down_isReady;
  wire                execute_ctrl5_down_LANE_SEL_lane0;
  wire       [63:0]   execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl5_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl5_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl4_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [63:0]   execute_ctrl4_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl3_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  wire       [63:0]   execute_ctrl3_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  wire       [4:0]    execute_ctrl4_down_RD_PHYS_lane1;
  wire                execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                execute_ctrl4_down_COMMIT_lane1;
  reg                 execute_ctrl4_up_RD_ENABLE_lane1;
  wire                execute_ctrl4_down_LANE_SEL_lane1;
  wire       [31:0]   execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  reg        [31:0]   execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire                execute_ctrl2_down_COMMIT_lane1;
  wire                execute_ctrl2_down_LANE_SEL_lane1;
  wire       [31:0]   execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  wire       [4:0]    execute_ctrl4_down_RD_PHYS_lane0;
  wire                execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [15:0]   execute_ctrl3_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl3_down_COMMIT_lane0;
  wire                execute_ctrl3_down_isReady;
  wire                execute_ctrl3_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire                execute_ctrl2_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  wire                FpuUnpackerPlugin_logic_unpacker_node_1_isValid;
  wire                FpuUnpackerPlugin_logic_unpacker_node_0_isValid;
  reg        [0:0]    FpuUnpackerPlugin_logic_unpacker_node_1_input_source;
  reg                 FpuUnpackerPlugin_logic_unpacker_node_2_valid;
  reg                 FpuUnpackerPlugin_logic_unpacker_node_1_valid;
  wire                execute_ctrl2_down_FpuUnpackerPlugin_SEL_I2F_lane0;
  wire                execute_ctrl2_down_FpuUnpack_RS3_badBoxing_HIT_lane0;
  wire       [0:0]    execute_ctrl2_down_RS3_RFID_lane0;
  reg                 execute_ctrl2_up_RS3_ENABLE_lane0;
  reg        [1:0]    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_sign;
  reg        [11:0]   execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mantissa;
  wire       [1:0]    execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_sign;
  reg        [10:0]   execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa;
  wire                execute_ctrl2_down_FpuUnpack_RS3_IS_SUBNORMAL_lane0;
  wire                execute_ctrl2_down_FpuUnpack_RS2_badBoxing_HIT_lane0;
  wire       [0:0]    execute_ctrl2_down_RS2_RFID_lane0;
  reg                 execute_ctrl2_up_RS2_ENABLE_lane0;
  reg        [1:0]    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign;
  reg        [11:0]   execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa;
  wire       [1:0]    execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_sign;
  reg        [10:0]   execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa;
  wire                execute_ctrl2_down_FpuUnpack_RS2_IS_SUBNORMAL_lane0;
  wire                execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0;
  wire       [0:0]    execute_ctrl2_down_RS1_RFID_lane0;
  reg                 execute_ctrl2_up_RS1_ENABLE_lane0;
  reg        [1:0]    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign;
  reg        [11:0]   execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa;
  wire       [1:0]    execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode;
  reg                 execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_quiet;
  reg                 execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_sign;
  reg        [10:0]   execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent;
  reg        [51:0]   execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa;
  wire       [0:0]    execute_ctrl2_down_FpuUtils_FORMAT_lane0;
  wire                execute_ctrl2_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1;
  wire                decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1;
  wire                decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  wire                decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  wire                decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  wire       [11:0]   decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [3:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [3:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [31:0]   decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0;
  wire                decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0;
  wire                decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0;
  wire                decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [11:0]   decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [3:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [3:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [31:0]   decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                decode_ctrls_1_up_isValid;
  reg                 decode_ctrls_1_down_ready;
  wire                execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
  wire                execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire                execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  wire                execute_ctrl7_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire                execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  wire                execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  wire                execute_ctrl3_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  wire                execute_ctrl9_down_BYPASSED_AT_10_lane0;
  reg        [0:0]    execute_ctrl9_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl9_up_RD_PHYS_lane0;
  reg                 execute_ctrl9_up_RD_ENABLE_lane0;
  wire                execute_ctrl8_down_BYPASSED_AT_9_lane0;
  reg        [0:0]    execute_ctrl8_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl8_up_RD_PHYS_lane0;
  reg                 execute_ctrl8_up_RD_ENABLE_lane0;
  wire                execute_ctrl7_down_BYPASSED_AT_8_lane0;
  reg        [0:0]    execute_ctrl7_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl7_up_RD_PHYS_lane0;
  reg                 execute_ctrl7_up_RD_ENABLE_lane0;
  wire                execute_ctrl6_down_BYPASSED_AT_7_lane0;
  reg        [0:0]    execute_ctrl6_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl6_up_RD_PHYS_lane0;
  reg                 execute_ctrl6_up_RD_ENABLE_lane0;
  wire                execute_ctrl5_down_BYPASSED_AT_6_lane0;
  reg        [0:0]    execute_ctrl5_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl5_up_RD_PHYS_lane0;
  reg                 execute_ctrl5_up_RD_ENABLE_lane0;
  wire                execute_ctrl4_down_BYPASSED_AT_5_lane0;
  reg        [0:0]    execute_ctrl4_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl4_up_RD_PHYS_lane0;
  reg                 execute_ctrl4_up_RD_ENABLE_lane0;
  wire                execute_ctrl3_down_BYPASSED_AT_4_lane0;
  reg        [0:0]    execute_ctrl3_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl3_up_RD_PHYS_lane0;
  reg                 execute_ctrl3_up_RD_ENABLE_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_3_lane1;
  reg        [0:0]    execute_ctrl2_up_RD_RFID_lane1;
  reg        [4:0]    execute_ctrl2_up_RD_PHYS_lane1;
  reg                 execute_ctrl2_up_RD_ENABLE_lane1;
  wire                execute_ctrl1_down_BYPASSED_AT_2_lane1;
  reg        [0:0]    execute_ctrl1_up_RD_RFID_lane1;
  reg        [4:0]    execute_ctrl1_up_RD_PHYS_lane1;
  reg                 execute_ctrl1_up_RD_ENABLE_lane1;
  wire                execute_ctrl2_down_BYPASSED_AT_3_lane0;
  reg        [0:0]    execute_ctrl2_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl2_up_RD_PHYS_lane0;
  reg                 execute_ctrl2_up_RD_ENABLE_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_2_lane0;
  reg        [0:0]    execute_ctrl1_up_RD_RFID_lane0;
  reg        [4:0]    execute_ctrl1_up_RD_PHYS_lane0;
  reg                 execute_ctrl1_up_RD_ENABLE_lane0;
  reg                 decode_ctrls_1_up_TRAP_1;
  reg                 decode_ctrls_1_TRAP_1_bypass;
  wire       [15:0]   decode_ctrls_1_down_Decode_UOP_ID_1;
  wire                decode_ctrls_1_down_TRAP_1;
  wire       [0:0]    decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [31:0]   decode_ctrls_1_down_PC_1;
  wire                decode_ctrls_1_down_Prediction_ALIGN_REDO_1;
  wire                decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1;
  reg                 decode_ctrls_1_up_LANE_SEL_1;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1;
  wire       [31:0]   decode_ctrls_1_down_Decode_UOP_1;
  wire                decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1;
  reg                 decode_ctrls_1_down_Decode_LEGAL_1;
  wire       [4:0]    decode_ctrls_1_down_RS3_PHYS_1;
  wire       [0:0]    decode_ctrls_1_down_RS3_RFID_1;
  wire                decode_ctrls_1_down_RS3_ENABLE_1;
  wire       [4:0]    decode_ctrls_1_down_RD_PHYS_1;
  wire       [0:0]    decode_ctrls_1_down_RD_RFID_1;
  reg                 decode_ctrls_1_down_RD_ENABLE_1;
  wire       [4:0]    decode_ctrls_1_down_RS2_PHYS_1;
  wire       [0:0]    decode_ctrls_1_down_RS2_RFID_1;
  wire                decode_ctrls_1_down_RS2_ENABLE_1;
  wire       [4:0]    decode_ctrls_1_down_RS1_PHYS_1;
  wire       [0:0]    decode_ctrls_1_down_RS1_RFID_1;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_1;
  wire                decode_ctrls_1_down_RS1_ENABLE_1;
  wire                decode_ctrls_1_lane1_upIsCancel;
  wire                decode_ctrls_1_lane1_downIsCancel;
  reg                 decode_ctrls_1_up_TRAP_0;
  reg                 decode_ctrls_1_TRAP_0_bypass;
  wire       [15:0]   decode_ctrls_1_down_Decode_UOP_ID_0;
  wire                decode_ctrls_1_up_isReady;
  wire                decode_ctrls_1_down_TRAP_0;
  wire       [0:0]    decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [31:0]   decode_ctrls_1_down_PC_0;
  wire                decode_ctrls_1_down_Prediction_ALIGN_REDO_0;
  wire                decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  reg                 decode_ctrls_1_up_LANE_SEL_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_UOP_0;
  wire                decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0;
  reg                 decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [4:0]    decode_ctrls_1_down_RS3_PHYS_0;
  wire       [0:0]    decode_ctrls_1_down_RS3_RFID_0;
  wire                decode_ctrls_1_down_RS3_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RD_PHYS_0;
  wire       [0:0]    decode_ctrls_1_down_RD_RFID_0;
  reg                 decode_ctrls_1_down_RD_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS2_PHYS_0;
  wire       [0:0]    decode_ctrls_1_down_RS2_RFID_0;
  wire                decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS1_PHYS_0;
  wire       [0:0]    decode_ctrls_1_down_RS1_RFID_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_1_down_RS1_ENABLE_0;
  wire                decode_ctrls_1_up_isCanceling;
  wire                decode_ctrls_1_up_ready;
  reg                 decode_ctrls_1_up_valid;
  wire                decode_ctrls_1_up_isMoving;
  wire                execute_ctrl2_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_COMPLETED_lane0;
  wire                execute_ctrl2_down_COMPLETED_lane0;
  wire                execute_ctrl2_COMPLETED_lane0_bypass;
  wire                execute_ctrl8_down_COMPLETION_AT_8_lane0;
  reg                 execute_ctrl8_up_COMPLETED_lane0;
  wire                execute_ctrl8_COMPLETED_lane0_bypass;
  wire                execute_ctrl5_down_COMPLETION_AT_5_lane0;
  reg                 execute_ctrl5_up_COMPLETED_lane0;
  wire                execute_ctrl5_COMPLETED_lane0_bypass;
  wire                execute_ctrl3_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_COMPLETED_lane0;
  wire                execute_ctrl3_down_COMPLETED_lane0;
  wire                execute_ctrl3_COMPLETED_lane0_bypass;
  wire                execute_ctrl11_down_COMPLETION_AT_11_lane0;
  reg                 execute_ctrl11_up_COMPLETED_lane0;
  wire                execute_ctrl11_COMPLETED_lane0_bypass;
  wire                execute_ctrl7_down_COMPLETION_AT_7_lane0;
  reg                 execute_ctrl7_up_COMPLETED_lane0;
  wire                execute_ctrl7_COMPLETED_lane0_bypass;
  wire                execute_ctrl4_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_COMPLETED_lane0;
  wire                execute_ctrl4_down_COMPLETED_lane0;
  wire                execute_ctrl4_COMPLETED_lane0_bypass;
  wire                execute_ctrl11_down_COMPLETED_lane0;
  wire                execute_ctrl10_down_COMPLETED_lane0;
  reg                 execute_ctrl10_up_LANE_SEL_lane0;
  wire                execute_ctrl9_down_COMPLETED_lane0;
  wire                execute_ctrl8_down_COMPLETED_lane0;
  wire                execute_ctrl7_down_COMPLETED_lane0;
  wire                execute_ctrl6_down_COMPLETED_lane0;
  wire                execute_ctrl5_down_COMPLETED_lane0;
  reg                 execute_ctrl1_up_LANE_SEL_lane0;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [31:0]   execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire                execute_ctrl4_down_early1_BranchPlugin_SEL_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1;
  wire       [15:0]   execute_ctrl4_down_Decode_UOP_ID_lane1;
  wire       [0:0]    execute_ctrl4_down_LANE_AGE_lane1;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_shifter_3;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_shifter_2;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [3:0]    execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [3:0]    execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [11:0]   execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [31:0]   execute_ctrl4_down_PC_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_SEL_lane1;
  wire                execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  wire       [31:0]   execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  wire       [31:0]   execute_ctrl4_down_Decode_UOP_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  wire       [1:0]    execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  wire       [31:0]   execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire       [31:0]   execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [31:0]   execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire                execute_ctrl4_down_early0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_shifter_3;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [3:0]    execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [3:0]    execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [11:0]   execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire       [31:0]   execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire       [1:0]    execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [31:0]   execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [31:0]   execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0;
  reg                 execute_ctrl11_up_COMMIT_lane0;
  reg                 execute_ctrl11_up_LANE_SEL_lane0;
  reg                 execute_ctrl8_up_COMMIT_lane0;
  reg                 execute_ctrl8_up_LANE_SEL_lane0;
  reg                 execute_ctrl5_up_COMMIT_lane0;
  reg                 execute_ctrl5_up_LANE_SEL_lane0;
  reg                 execute_ctrl7_up_COMMIT_lane0;
  reg                 execute_ctrl7_up_LANE_SEL_lane0;
  reg                 execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  reg                 execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  reg                 execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  reg                 execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  reg                 execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  wire                execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  wire                execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  wire                execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  wire                execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  wire                execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  wire                execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX;
  wire                execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_UF;
  wire                execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_OF;
  wire                execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_DZ;
  wire                execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NV;
  wire                execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  wire                execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  wire                execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  wire                execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  wire                execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  wire                execute_ctrl4_down_COMPLETION_AT_4_lane1;
  reg                 execute_ctrl4_up_COMPLETED_lane1;
  wire                execute_ctrl4_down_COMPLETED_lane1;
  wire                execute_ctrl4_COMPLETED_lane1_bypass;
  wire                execute_ctrl2_down_COMPLETION_AT_2_lane1;
  reg                 execute_ctrl2_up_COMPLETED_lane1;
  wire                execute_ctrl2_down_COMPLETED_lane1;
  wire                execute_ctrl2_COMPLETED_lane1_bypass;
  reg                 execute_ctrl3_up_LANE_SEL_lane1;
  reg                 execute_ctrl1_up_LANE_SEL_lane1;
  wire                PrefetcherRptPlugin_logic_pip_node_2_isReady;
  wire                PrefetcherRptPlugin_logic_pip_node_2_isValid;
  wire                PrefetcherRptPlugin_logic_pip_node_0_isReady;
  wire                PrefetcherRptPlugin_logic_pip_node_1_isValid;
  wire                PrefetcherRptPlugin_logic_pip_node_0_isValid;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_valid;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_valid;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_TAG_HIT;
  wire                PrefetcherRptPlugin_logic_pip_node_2_isFiring;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_NEW_BLOCK;
  reg        [31:0]   PrefetcherRptPlugin_logic_pip_node_2_PROBE_pc;
  reg        [31:0]   PrefetcherRptPlugin_logic_pip_node_2_PROBE_address;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_load;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_store;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_trap;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_io;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_prefetchFailed;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_PROBE_miss;
  wire       [11:0]   PrefetcherRptPlugin_logic_pip_node_2_STRIDE;
  reg        [14:0]   PrefetcherRptPlugin_logic_pip_node_2_ENTRY_tag;
  reg        [15:0]   PrefetcherRptPlugin_logic_pip_node_2_ENTRY_address;
  reg        [11:0]   PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride;
  reg        [4:0]    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score;
  reg        [2:0]    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_advance;
  reg                 PrefetcherRptPlugin_logic_pip_node_2_ENTRY_missed;
  reg        [15:0]   PrefetcherRptPlugin_logic_pip_node_2_STRIDE_EXTENDED;
  wire                PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT;
  wire                PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK;
  wire       [15:0]   PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED;
  wire                PrefetcherRptPlugin_logic_pip_node_1_TAG_HIT;
  reg        [31:0]   PrefetcherRptPlugin_logic_pip_node_1_PROBE_pc;
  reg        [31:0]   PrefetcherRptPlugin_logic_pip_node_1_PROBE_address;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_load;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_store;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_trap;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_io;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_prefetchFailed;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_PROBE_miss;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_valid;
  reg        [6:0]    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_address;
  reg        [14:0]   PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_tag;
  reg        [15:0]   PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_address;
  reg        [11:0]   PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_stride;
  reg        [4:0]    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_score;
  reg        [2:0]    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_advance;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_missed;
  reg        [14:0]   PrefetcherRptPlugin_logic_pip_node_1_ENTRY_tag;
  reg        [15:0]   PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address;
  reg        [11:0]   PrefetcherRptPlugin_logic_pip_node_1_ENTRY_stride;
  reg        [4:0]    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_score;
  reg        [2:0]    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_advance;
  reg                 PrefetcherRptPlugin_logic_pip_node_1_ENTRY_missed;
  wire                PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_valid;
  wire       [6:0]    PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_address;
  wire       [14:0]   PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_tag;
  wire       [15:0]   PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_address;
  wire       [11:0]   PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_stride;
  wire       [4:0]    PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_score;
  wire       [2:0]    PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_advance;
  wire                PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_missed;
  wire                PrefetcherRptPlugin_logic_pip_node_0_isFiring;
  wire       [31:0]   PrefetcherRptPlugin_logic_pip_node_0_PROBE_pc;
  wire       [31:0]   PrefetcherRptPlugin_logic_pip_node_0_PROBE_address;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_load;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_store;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_trap;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_io;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_prefetchFailed;
  wire                PrefetcherRptPlugin_logic_pip_node_0_PROBE_miss;
  wire                PrefetcherRptPlugin_logic_pip_node_0_valid;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1;
  wire       [15:0]   execute_ctrl2_down_Decode_UOP_ID_lane1;
  wire       [0:0]    execute_ctrl2_down_LANE_AGE_lane1;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_shifter_3;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_shifter_2;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [3:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [3:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [11:0]   execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
  wire                execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  wire       [31:0]   execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_3;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [3:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [3:0]    execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [11:0]   execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [31:0]   execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire                FpuPackerPlugin_logic_pip_node_1_isReady;
  wire                FpuPackerPlugin_logic_pip_node_0_isValid;
  wire                FpuPackerPlugin_logic_pip_node_0_isReady;
  reg        [4:0]    FpuPackerPlugin_logic_pip_node_1_s0_GROUP_OH;
  reg        [15:0]   FpuPackerPlugin_logic_pip_node_1_Decode_UOP_ID;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NX;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_UF;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_OF;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_DZ;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NV;
  reg                 FpuPackerPlugin_logic_pip_node_1_valid;
  wire                FpuPackerPlugin_logic_pip_node_0_ready;
  wire                FpuPackerPlugin_logic_pip_node_1_ready;
  wire                FpuPackerPlugin_logic_pip_node_2_ready;
  reg        [51:0]   FpuPackerPlugin_logic_pip_node_2_s1_MAN_RESULT;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NX;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_UF;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_OF;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_DZ;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NV;
  reg        [15:0]   FpuPackerPlugin_logic_pip_node_2_Decode_UOP_ID;
  reg                 FpuPackerPlugin_logic_pip_node_2_valid;
  reg        [4:0]    FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH;
  reg                 FpuPackerPlugin_logic_pip_node_2_s1_ROUNDING_INCR;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_subnormal_ENABLE;
  reg        [1:0]    FpuPackerPlugin_logic_pip_node_2_s1_roundAdjusted;
  reg                 FpuPackerPlugin_logic_pip_node_2_s1_manLsb;
  reg        [2:0]    FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE;
  reg        [1:0]    FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_VALUE_quiet;
  reg                 FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign;
  reg        [12:0]   FpuPackerPlugin_logic_pip_node_2_s0_VALUE_exponent;
  reg        [53:0]   FpuPackerPlugin_logic_s2_mr;
  wire                FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW;
  wire                FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW;
  wire       [11:0]   FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN;
  wire       [10:0]   FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX;
  reg        [0:0]    FpuPackerPlugin_logic_pip_node_2_s0_FORMAT;
  wire       [12:0]   FpuPackerPlugin_logic_pip_node_2_s2_EXP;
  wire                FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL;
  reg        [12:0]   FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  reg        [10:0]   FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL;
  wire       [51:0]   FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT;
  wire       [12:0]   FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT;
  wire       [12:0]   FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR;
  wire                FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR;
  reg        [2:0]    FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE;
  wire                FpuPackerPlugin_logic_pip_node_1_s1_manLsb;
  wire       [1:0]    FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted;
  reg        [0:0]    FpuPackerPlugin_logic_pip_node_1_s0_FORMAT;
  wire                FpuPackerPlugin_logic_pip_node_1_isValid;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_subnormal_ENABLE;
  reg        [54:0]   _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter;
  reg        [54:0]   _zz_when_Utils_l1585_3;
  reg        [54:0]   _zz_when_Utils_l1585_4;
  reg        [54:0]   _zz_when_Utils_l1585_5;
  reg        [54:0]   _zz_when_Utils_l1585_6;
  reg        [54:0]   _zz_when_Utils_l1585_7;
  wire       [12:0]   FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE;
  reg        [10:0]   FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL;
  reg        [53:0]   FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED;
  reg        [1:0]    FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_VALUE_quiet;
  reg                 FpuPackerPlugin_logic_pip_node_1_s0_VALUE_sign;
  reg        [12:0]   FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  reg        [53:0]   FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mantissa;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE;
  wire       [10:0]   FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL;
  reg        [4:0]    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH;
  wire                FpuPackerPlugin_logic_pip_node_0_valid;
  wire       [15:0]   FpuPackerPlugin_logic_pip_node_0_Decode_UOP_ID;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_UF;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_OF;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_DZ;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NV;
  wire       [2:0]    FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE;
  wire       [0:0]    FpuPackerPlugin_logic_pip_node_0_s0_FORMAT;
  wire       [1:0]    FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet;
  wire                FpuPackerPlugin_logic_pip_node_0_s0_VALUE_sign;
  wire       [12:0]   FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_1_isReady;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_1_isValid;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_0_isValid;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_0_isReady;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_ops_pip_node_1_SB_PTR;
  reg                 LsuPlugin_logic_storeBuffer_ops_pip_node_2_valid;
  reg                 LsuPlugin_logic_storeBuffer_ops_pip_node_1_valid;
  reg                 LsuPlugin_logic_storeBuffer_ops_pip_node_0_ready;
  reg                 LsuPlugin_logic_storeBuffer_ops_pip_node_1_ready;
  wire       [1:0]    execute_ctrl4_down_AguPlugin_SIZE_lane0;
  wire       [31:0]   execute_ctrl4_down_PC_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  wire                execute_ctrl4_down_LANE_SEL_lane0;
  reg                 execute_ctrl4_up_COMMIT_lane0;
  reg                 execute_ctrl4_COMMIT_lane0_bypass;
  reg                 execute_ctrl4_up_TRAP_lane0;
  wire                execute_ctrl4_down_TRAP_lane0;
  reg                 execute_ctrl4_TRAP_lane0_bypass;
  wire                execute_ctrl4_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0;
  wire       [11:0]   execute_ctrl4_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  wire                execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0;
  wire                execute_ctrl4_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire                execute_ctrl4_down_MMU_HAZARD_lane0;
  wire                execute_ctrl4_down_MMU_REFILL_lane0;
  wire                execute_ctrl4_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire       [0:0]    execute_ctrl4_down_LANE_AGE_lane0;
  wire       [5:0]    execute_ctrl4_down_LsuPlugin_SB_PTR_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire       [31:0]   execute_ctrl4_down_integer_RS2_lane0;
  wire       [31:0]   execute_ctrl4_down_Decode_UOP_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  wire       [15:0]   execute_ctrl4_down_Decode_UOP_ID_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  reg        [63:0]   execute_ctrl4_up_float_RS2_lane0;
  wire                execute_ctrl4_down_AguPlugin_FLOAT_lane0;
  reg        [31:0]   execute_ctrl4_up_integer_RS2_lane0;
  wire                execute_ctrl3_down_MMU_HAZARD_lane0;
  wire                execute_ctrl3_down_MMU_REFILL_lane0;
  wire                execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  wire                execute_ctrl3_down_MMU_ALLOW_READ_lane0;
  wire                execute_ctrl3_down_MMU_ALLOW_WRITE_lane0;
  wire                execute_ctrl3_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl3_down_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire                execute_ctrl3_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg                 execute_ctrl4_LsuL1_SEL_lane0_bypass;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl4_up_LsuL1_SEL_lane0;
  reg                 execute_ctrl3_LsuL1_SEL_lane0_bypass;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl3_up_LsuL1_SEL_lane0;
  wire       [31:0]   execute_ctrl3_down_MMU_TRANSLATED_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  wire       [63:0]   execute_ctrl2_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  wire       [5:0]    execute_ctrl2_down_LsuPlugin_SB_PTR_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
  wire       [11:0]   execute_ctrl2_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl2_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl2_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl2_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl2_down_LsuL1_STORE_lane0;
  wire                execute_ctrl2_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl2_down_LsuL1_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_LsuL1_SIZE_lane0;
  wire       [7:0]    execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                execute_ctrl2_down_LsuL1_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl2_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl2_down_AguPlugin_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl2_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire       [1:0]    execute_ctrl3_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl3_down_LsuL1_STORE_lane0;
  wire                execute_ctrl3_down_LsuL1_LOAD_lane0;
  wire                execute_ctrl3_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl3_down_LsuL1_SEL_lane0;
  reg                 _zz_2;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_ops_pip_node_2_SB_PTR;
  reg        [31:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_address;
  reg        [63:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_data;
  reg        [1:0]    LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_size;
  reg        [11:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_storeId;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_2_ready;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_2_isValid;
  wire       [31:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address;
  wire       [63:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_data;
  wire       [1:0]    LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_size;
  wire       [11:0]   LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_storeId;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_0_isFiring;
  wire       [5:0]    LsuPlugin_logic_storeBuffer_ops_pip_node_0_SB_PTR;
  wire                LsuPlugin_logic_storeBuffer_ops_pip_node_0_valid;
  wire       [31:0]   execute_ctrl0_down_Decode_UOP_lane0;
  wire                execute_ctrl4_down_FpuCsrPlugin_DIRTY_lane0;
  wire                execute_ctrl4_down_COMMIT_lane0;
  wire                execute_ctrl4_down_isReady;
  wire       [2:0]    execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  wire       [31:0]   fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
  wire       [3:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
  wire       [3:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3;
  wire       [9:0]    fetch_logic_ctrls_2_down_Fetch_ID;
  wire                fetch_logic_ctrls_2_down_isCancel;
  wire                fetch_logic_ctrls_2_down_ready;
  wire                decode_ctrls_0_up_isCancel;
  wire                fetch_logic_ctrls_2_down_valid;
  wire                fetch_logic_ctrls_2_down_isValid;
  wire                decode_ctrls_0_up_valid;
  wire                decode_ctrls_0_up_Prediction_ALIGN_REDO_1;
  wire       [3:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [3:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [31:0]   decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1;
  wire                decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1;
  wire                decode_ctrls_0_up_TRAP_1;
  wire       [1:0]    decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1;
  wire                decode_ctrls_0_up_Prediction_WORD_JUMPED_1;
  wire       [31:0]   decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1;
  wire       [3:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1;
  wire       [3:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1;
  wire       [11:0]   decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [9:0]    decode_ctrls_0_up_Fetch_ID_1;
  wire       [9:0]    decode_ctrls_0_up_Decode_DOP_ID_1;
  wire       [31:0]   decode_ctrls_0_up_PC_1;
  wire       [0:0]    decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1;
  reg                 decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_1;
  wire                decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  wire       [3:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [3:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  wire                decode_ctrls_0_up_TRAP_0;
  wire       [1:0]    decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0;
  wire                decode_ctrls_0_up_Prediction_WORD_JUMPED_0;
  wire       [31:0]   decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  wire       [3:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  wire       [3:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  wire       [11:0]   decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [9:0]    decode_ctrls_0_up_Fetch_ID_0;
  wire       [9:0]    decode_ctrls_0_up_Decode_DOP_ID_0;
  wire       [31:0]   decode_ctrls_0_up_PC_0;
  wire       [0:0]    decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  reg                 decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_up_isFiring;
  wire       [3:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
  wire       [1:0]    fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
  wire       [3:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [31:0]   execute_ctrl2_down_PC_lane1;
  wire       [1:0]    execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire       [31:0]   execute_ctrl2_down_Decode_UOP_lane1;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [1:0]    execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl2_up_COMMIT_lane0;
  wire                execute_ctrl2_down_COMMIT_lane0;
  reg                 execute_ctrl2_COMMIT_lane0_bypass;
  reg                 execute_ctrl2_up_TRAP_lane0;
  wire                execute_ctrl2_down_TRAP_lane0;
  reg                 execute_ctrl2_TRAP_lane0_bypass;
  wire                execute_ctrl2_down_early0_EnvPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_Decode_UOP_lane0;
  wire       [31:0]   execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
  wire                execute_ctrl2_down_DivPlugin_REM_lane0;
  wire                execute_ctrl4_down_MulPlugin_HIGH_lane0;
  wire                execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  wire       [110:0]  execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  wire       [5:0]    execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  wire       [46:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [63:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [5:0]    execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [22:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [22:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [39:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [39:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [56:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [56:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [5:0]    execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  wire       [46:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [63:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [5:0]    execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [22:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [22:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [39:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [39:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [56:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [56:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [5:0]    execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  wire       [22:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  wire       [22:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  wire       [39:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  wire       [39:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  wire       [56:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  wire       [56:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg        [53:0]   execute_ctrl2_down_MUL_SRC2_lane0;
  reg        [53:0]   execute_ctrl2_down_MUL_SRC1_lane0;
  wire                execute_ctrl2_down_isReady;
  reg        [63:0]   execute_ctrl2_up_float_RS3_lane0;
  reg        [63:0]   execute_ctrl2_up_float_RS2_lane0;
  reg        [63:0]   execute_ctrl2_up_float_RS1_lane0;
  reg        [0:0]    FpuUnpackerPlugin_logic_unpacker_node_2_input_source;
  wire                FpuUnpackerPlugin_logic_unpacker_node_2_isValid;
  reg        [5:0]    FpuUnpackerPlugin_logic_unpacker_node_2_setup_shiftBy;
  reg        [51:0]   FpuUnpackerPlugin_logic_unpacker_node_2_input_args_data;
  wire       [5:0]    FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy;
  reg        [51:0]   FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data;
  wire       [0:0]    FpuUnpackerPlugin_logic_unpacker_node_0_input_source;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_node_0_input_args_data;
  wire                FpuUnpackerPlugin_logic_unpacker_node_0_valid;
  wire                FpuAddSharedPlugin_logic_pip_node_3_isValid;
  wire                FpuAddSharedPlugin_logic_pip_node_3_isReady;
  wire                FpuAddSharedPlugin_logic_pip_node_2_isValid;
  wire                FpuAddSharedPlugin_logic_pip_node_2_isReady;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_adder_math_roundingScrap;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xySign;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_3_inserter_GROUP_OH;
  reg        [15:0]   FpuAddSharedPlugin_logic_pip_node_3_Decode_UOP_ID;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NX;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_UF;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_OF;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_DZ;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NV;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_RDN;
  reg        [2:0]    FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE;
  reg        [0:0]    FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT;
  wire                FpuAddSharedPlugin_logic_pip_node_1_isValid;
  wire                FpuAddSharedPlugin_logic_pip_node_1_isReady;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xySign;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_2_inserter_GROUP_OH;
  reg        [15:0]   FpuAddSharedPlugin_logic_pip_node_2_Decode_UOP_ID;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NX;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_UF;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_OF;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_DZ;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NV;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_RDN;
  reg        [2:0]    FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE;
  reg        [0:0]    FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT;
  wire                FpuAddSharedPlugin_logic_pip_node_0_isReady;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_passThrough;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_needSub;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_1_inserter_GROUP_OH;
  reg        [15:0]   FpuAddSharedPlugin_logic_pip_node_1_Decode_UOP_ID;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NX;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_UF;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_OF;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_DZ;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NV;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_RDN;
  reg        [2:0]    FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE;
  reg        [0:0]    FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_valid;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_valid;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_valid;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_valid;
  wire                FpuAddSharedPlugin_logic_pip_node_0_ready;
  wire                FpuAddSharedPlugin_logic_pip_node_1_ready;
  wire                FpuAddSharedPlugin_logic_pip_node_2_ready;
  wire                FpuAddSharedPlugin_logic_pip_node_3_ready;
  wire                FpuAddSharedPlugin_logic_pip_node_4_ready;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NX;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_UF;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_OF;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_DZ;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NV;
  reg        [15:0]   FpuAddSharedPlugin_logic_pip_node_4_Decode_UOP_ID;
  reg        [2:0]    FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE;
  reg        [0:0]    FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT;
  reg                 execute_ctrl9_up_LANE_SEL_lane0;
  reg                 execute_ctrl6_up_LANE_SEL_lane0;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_4_inserter_GROUP_OH;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_RDN;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_norm_xyMantissaZero;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceZero;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceInfinity;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceNan;
  wire                FpuAddSharedPlugin_logic_pip_node_4_adder_result_NV;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_sign;
  reg        [11:0]   FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_exponent;
  reg        [51:0]   FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mantissa;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_sign;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_exponent;
  reg        [104:0]  FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mantissa;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_norm_infinityNan;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_math_roundingScrap;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xySign;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_sign;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_4_adder_result_mantissa;
  reg        [107:0]  FpuAddSharedPlugin_logic_pip_node_4_adder_math_xyMantissa;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent;
  reg        [6:0]    FpuAddSharedPlugin_logic_pip_node_4_adder_norm_shift;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent;
  wire                FpuAddSharedPlugin_logic_pip_node_3_adder_norm_xyMantissaZero;
  wire                FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceNan;
  wire                FpuAddSharedPlugin_logic_pip_node_3_adder_norm_infinityNan;
  wire                FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceZero;
  wire                FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceInfinity;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_sign;
  reg        [11:0]   FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent;
  reg        [51:0]   FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mantissa;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_sign;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent;
  reg        [104:0]  FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mantissa;
  wire       [6:0]    FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh;
  reg        [107:0]  FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa;
  reg        [105:0]  FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xMantissa;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_needSub;
  reg        [106:0]  FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_yMantissa;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_sign;
  reg        [11:0]   FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent;
  reg        [51:0]   FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mantissa;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_sign;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent;
  reg        [104:0]  FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mantissa;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_adder_math_roundingScrap;
  reg                 FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_passThrough;
  reg        [107:0]  FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_shifter;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent;
  wire       [106:0]  FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissa;
  wire       [107:0]  FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter;
  reg        [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter;
  reg        [107:0]  _zz_when_Utils_l1585_8;
  reg        [107:0]  _zz_when_Utils_l1585_9;
  reg        [107:0]  _zz_when_Utils_l1585_10;
  reg        [107:0]  _zz_when_Utils_l1585_11;
  reg        [107:0]  _zz_when_Utils_l1585_12;
  reg        [107:0]  _zz_when_Utils_l1585_13;
  reg        [6:0]    FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat;
  wire       [105:0]  FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted;
  wire       [105:0]  FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa;
  wire                FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xySign;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_sign;
  reg        [11:0]   FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent;
  reg        [51:0]   FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mantissa;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_quiet;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_sign;
  reg        [12:0]   FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent;
  reg        [104:0]  FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mantissa;
  reg                 FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger;
  wire       [6:0]    FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_passThrough;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_needSub;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_absRs1Bigger;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual;
  wire                FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentBigger;
  wire       [11:0]   FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21;
  reg        [1:0]    FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH;
  wire                FpuAddSharedPlugin_logic_pip_node_0_isValid;
  wire                FpuAddSharedPlugin_logic_pip_node_0_valid;
  wire       [15:0]   FpuAddSharedPlugin_logic_pip_node_0_Decode_UOP_ID;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_UF;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_OF;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_DZ;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NV;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_RDN;
  wire       [2:0]    FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE;
  wire       [0:0]    FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT;
  wire       [1:0]    FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_sign;
  wire       [11:0]   FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  wire       [51:0]   FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa;
  wire       [1:0]    FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet;
  wire                FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_sign;
  wire       [12:0]   FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  wire       [104:0]  FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa;
  wire                execute_ctrl4_down_SrcStageables_UNSIGNED_lane1;
  wire                execute_ctrl4_down_SrcStageables_ZERO_lane1;
  wire                execute_ctrl4_down_SrcStageables_REVERT_lane1;
  wire       [31:0]   execute_ctrl3_down_PC_lane1;
  wire       [31:0]   execute_ctrl3_down_integer_RS2_lane1;
  wire       [1:0]    execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [31:0]   execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   execute_ctrl3_down_integer_RS1_lane1;
  wire       [0:0]    execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [31:0]   execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  wire       [31:0]   execute_ctrl3_down_Decode_UOP_lane1;
  reg                 execute_ctrl4_up_LANE_SEL_lane1;
  reg                 execute_ctrl2_up_LANE_SEL_lane1;
  wire                execute_ctrl2_down_SrcStageables_UNSIGNED_lane1;
  wire                execute_ctrl2_down_SrcStageables_ZERO_lane1;
  wire                execute_ctrl2_down_SrcStageables_REVERT_lane1;
  wire       [31:0]   execute_ctrl1_down_PC_lane1;
  wire       [31:0]   execute_ctrl1_down_integer_RS2_lane1;
  wire       [1:0]    execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [31:0]   execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   execute_ctrl1_down_integer_RS1_lane1;
  wire       [0:0]    execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [31:0]   execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  wire       [31:0]   execute_ctrl1_down_Decode_UOP_lane1;
  wire                execute_ctrl4_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl4_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl4_down_SrcStageables_REVERT_lane0;
  wire       [31:0]   execute_ctrl3_down_PC_lane0;
  wire       [31:0]   execute_ctrl3_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [31:0]   execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl3_down_integer_RS1_lane0;
  wire       [0:0]    execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [31:0]   execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  wire       [31:0]   execute_ctrl3_down_Decode_UOP_lane0;
  reg                 execute_ctrl3_up_LANE_SEL_lane0;
  wire       [1:0]    execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl4_up_LANE_SEL_lane0;
  reg                 execute_ctrl2_up_LANE_SEL_lane0;
  wire                execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl2_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl2_down_SrcStageables_REVERT_lane0;
  wire       [31:0]   execute_ctrl1_down_PC_lane0;
  wire       [31:0]   execute_ctrl1_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [31:0]   execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl1_down_integer_RS1_lane0;
  wire       [0:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [31:0]   execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  wire       [31:0]   execute_ctrl1_down_Decode_UOP_lane0;
  wire       [2:0]    execute_ctrl2_down_early0_EnvPlugin_OP_lane0;
  wire       [31:0]   execute_ctrl2_down_PC_lane0;
  wire       [0:0]    execute_ctrl2_down_LANE_AGE_lane0;
  wire       [15:0]   execute_ctrl2_down_Decode_UOP_ID_lane0;
  wire                decode_ctrls_1_lane0_upIsCancel;
  wire                decode_ctrls_1_lane0_downIsCancel;
  wire       [9:0]    decode_ctrls_0_down_Decode_DOP_ID_1;
  wire       [9:0]    decode_ctrls_0_down_Fetch_ID_1;
  wire       [31:0]   decode_ctrls_0_down_PC_1;
  wire                decode_ctrls_0_up_LANE_SEL_1;
  wire                decode_ctrls_0_lane1_upIsCancel;
  wire                decode_ctrls_0_lane1_downIsCancel;
  wire       [9:0]    decode_ctrls_0_down_Decode_DOP_ID_0;
  wire       [9:0]    decode_ctrls_0_down_Fetch_ID_0;
  wire       [31:0]   decode_ctrls_0_down_PC_0;
  wire                decode_ctrls_0_up_isReady;
  wire                decode_ctrls_0_up_LANE_SEL_0;
  wire                decode_ctrls_0_lane0_upIsCancel;
  wire                decode_ctrls_0_lane0_downIsCancel;
  wire       [9:0]    fetch_logic_ctrls_0_down_Fetch_ID;
  reg                 _zz_3;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire                fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_0_down_isReady;
  wire                fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3;
  wire       [11:0]   fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  reg                 _zz_4;
  wire       [1:0]    execute_ctrl0_down_AguPlugin_SIZE_lane0;
  wire                fetch_logic_ctrls_2_up_isCanceling;
  wire                fetch_logic_ctrls_2_down_isReady;
  wire                fetch_logic_ctrls_2_down_TRAP;
  wire                fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_2_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_HAZARD;
  wire                fetch_logic_ctrls_2_down_MMU_REFILL;
  wire                fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE;
  wire                fetch_logic_ctrls_2_down_MMU_PAGE_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_2_up_isCancel;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  wire       [31:0]   fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_2_up_isReady;
  wire                fetch_logic_ctrls_2_up_isValid;
  wire       [0:0]    fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [31:0]   fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_TRANSLATED;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [5:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
  wire       [63:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [63:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [63:0]   fetch_logic_ctrls_2_down_Fetch_WORD;
  wire       [31:0]   fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg        [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [5:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire       [0:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 fetch_logic_ctrls_1_up_valid;
  wire                fetch_logic_ctrls_1_up_ready;
  wire       [31:0]   fetch_logic_ctrls_0_down_Fetch_WORD_PC;
  reg                 _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
  reg                 _zz_5;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg                 _zz_6;
  wire       [255:0]  fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0;
  wire       [255:0]  fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1;
  reg                 _zz_7;
  wire                fetch_logic_ctrls_0_down_isFiring;
  reg        [31:0]   execute_ctrl4_up_integer_RS1_lane0;
  wire                execute_ctrl4_down_FpuMvPlugin_SEL_FLOAT_lane0;
  reg        [63:0]   execute_ctrl3_up_float_RS1_lane0;
  wire                execute_ctrl3_down_FpuMvPlugin_SEL_INT_lane0;
  wire                execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  wire                execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1;
  wire                execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1;
  wire                execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
  wire                execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1;
  wire       [1:0]    execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  wire                execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1;
  wire                execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1;
  wire                execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire                execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
  wire                execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1;
  wire       [1:0]    execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0;
  wire                execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
  wire                execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0;
  reg        [31:0]   execute_ctrl2_up_integer_RS2_lane0;
  reg        [31:0]   execute_ctrl2_up_integer_RS1_lane0;
  reg                 _zz_8;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_isValid;
  reg                 PrefetcherRptPlugin_logic_pip2_node_1_valid;
  reg                 PrefetcherRptPlugin_logic_pip2_node_0_ready;
  wire                PrefetcherRptPlugin_logic_pip2_node_1_ready;
  wire                PrefetcherRptPlugin_logic_pip2_node_1_isValid;
  wire       [31:0]   PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR;
  reg        [15:0]   PrefetcherRptPlugin_logic_pip2_node_1_MUL;
  reg        [31:0]   PrefetcherRptPlugin_logic_pip2_node_1_CMD_address;
  reg                 PrefetcherRptPlugin_logic_pip2_node_1_CMD_unique;
  reg        [2:0]    PrefetcherRptPlugin_logic_pip2_node_1_CMD_from;
  reg        [2:0]    PrefetcherRptPlugin_logic_pip2_node_1_CMD_to;
  reg        [11:0]   PrefetcherRptPlugin_logic_pip2_node_1_CMD_stride;
  wire       [15:0]   PrefetcherRptPlugin_logic_pip2_node_0_MUL;
  wire       [31:0]   PrefetcherRptPlugin_logic_pip2_node_0_CMD_address;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_CMD_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_pip2_node_0_CMD_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_pip2_node_0_CMD_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_pip2_node_0_CMD_stride;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_isFiring;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_isCancel;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_isReady;
  wire                PrefetcherRptPlugin_logic_pip2_node_0_valid;
  wire       [63:0]   execute_ctrl4_down_LsuL1_READ_DATA_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [7:0]    execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [7:0]    execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  wire       [7:0]    execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [63:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0;
  wire       [7:0]    execute_ctrl4_down_LsuL1_MASK_lane0;
  reg        [63:0]   execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
  wire                execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0;
  wire                execute_ctrl4_down_LsuL1_SEL_lane0;
  wire                execute_ctrl4_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl4_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl4_down_LsuL1_REFILL_HIT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1_FAULT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire                execute_ctrl4_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuL1_LOAD_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  wire       [0:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire                execute_ctrl4_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl4_down_LsuL1_STORE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  wire       [1:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [63:0]   execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [255:0]  execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0;
  wire       [255:0]  execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1;
  reg        [1:0]    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
  reg                 _zz_9;
  reg                 _zz_10;
  wire                execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                AlignerPlugin_api_singleFetch;
  wire                AlignerPlugin_api_downMoving;
  wire                AlignerPlugin_api_haltIt;
  reg                 DispatchPlugin_api_haltDispatch;
  wire                execute_freeze_valid;
  wire       [0:0]    execute_lane0_api_hartsInflight;
  wire                execute_lane0_ctrls_2_upIsCancel;
  wire                execute_lane0_ctrls_2_downIsCancel;
  wire                PrefetcherRptPlugin_io_valid;
  wire                PrefetcherRptPlugin_io_ready;
  wire       [31:0]   PrefetcherRptPlugin_io_payload_address;
  wire                PrefetcherRptPlugin_io_payload_unique;
  wire                CsrRamPlugin_api_holdRead;
  wire                CsrRamPlugin_api_holdWrite;
  reg                 CsrAccessPlugin_bus_decode_exception;
  wire                CsrAccessPlugin_bus_decode_read;
  wire                CsrAccessPlugin_bus_decode_write;
  wire       [11:0]   CsrAccessPlugin_bus_decode_address;
  reg                 CsrAccessPlugin_bus_decode_trap;
  wire                PrivilegedPlugin_api_lsuTriggerBus_load;
  wire                PrivilegedPlugin_api_lsuTriggerBus_store;
  wire       [31:0]   PrivilegedPlugin_api_lsuTriggerBus_virtual;
  wire       [1:0]    PrivilegedPlugin_api_lsuTriggerBus_size;
  wire                PrivilegedPlugin_api_harts_0_allowInterrupts;
  wire                PrivilegedPlugin_api_harts_0_allowException;
  wire                PrivilegedPlugin_api_harts_0_allowEbreakException;
  reg                 PrivilegedPlugin_api_harts_0_fpuEnable;
  reg                 TrapPlugin_api_harts_0_redo;
  reg                 TrapPlugin_api_harts_0_askWake;
  reg                 TrapPlugin_api_harts_0_rvTrap;
  wire                TrapPlugin_api_harts_0_fsmBusy;
  wire       [0:0]    execute_lane1_api_hartsInflight;
  wire                execute_lane1_ctrls_2_upIsCancel;
  wire                execute_lane1_ctrls_2_downIsCancel;
  reg        [2:0]    FpuCsrPlugin_api_rm;
  reg                 FpuCsrPlugin_api_flags_NX;
  reg                 FpuCsrPlugin_api_flags_UF;
  reg                 FpuCsrPlugin_api_flags_OF;
  reg                 FpuCsrPlugin_api_flags_DZ;
  reg                 FpuCsrPlugin_api_flags_NV;
  reg                 FpuCsrPlugin_api_gotDirty;
  wire                BtbPlugin_logic_pcPort_valid;
  wire                BtbPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   BtbPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid;
  wire                BtbPlugin_logic_historyPort_valid;
  wire       [11:0]   BtbPlugin_logic_historyPort_payload_history;
  wire                BtbPlugin_logic_flushPort_valid;
  wire                BtbPlugin_logic_flushPort_payload_self;
  wire                FetchL1Plugin_logic_bus_cmd_valid;
  wire                FetchL1Plugin_logic_bus_cmd_ready;
  wire       [0:0]    FetchL1Plugin_logic_bus_cmd_payload_id;
  wire       [31:0]   FetchL1Plugin_logic_bus_cmd_payload_address;
  wire                FetchL1Plugin_logic_bus_cmd_payload_io;
  wire                FetchL1Plugin_logic_bus_rsp_valid;
  wire                FetchL1Plugin_logic_bus_rsp_ready;
  wire       [0:0]    FetchL1Plugin_logic_bus_rsp_payload_id;
  wire       [255:0]  FetchL1Plugin_logic_bus_rsp_payload_data;
  wire                FetchL1Plugin_logic_bus_rsp_payload_error;
  reg                 FetchL1Plugin_logic_trapPort_valid;
  reg                 FetchL1Plugin_logic_trapPort_payload_exception;
  wire       [31:0]   FetchL1Plugin_logic_trapPort_payload_tval;
  wire       [0:0]    decode_logic_trapPending;
  wire       [0:0]    DispatchPlugin_logic_trapPendings;
  wire       [0:0]    execute_lane0_logic_trapPending;
  wire                early0_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   early0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   early0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   early0_IntAluPlugin_logic_alu_result;
  wire                early0_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_patched;
  wire                early0_BranchPlugin_logic_wb_valid;
  wire       [31:0]   early0_BranchPlugin_logic_wb_payload;
  wire                early0_BranchPlugin_logic_pcPort_valid;
  wire                early0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   early0_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    early0_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid;
  wire                early0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early0_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    early0_BranchPlugin_logic_historyPort_payload_age;
  wire                early0_BranchPlugin_logic_flushPort_valid;
  wire                LsuPlugin_logic_fpwb_valid;
  reg        [63:0]   LsuPlugin_logic_fpwb_payload;
  reg                 LsuPlugin_logic_trapPort_valid;
  reg                 LsuPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   LsuPlugin_logic_trapPort_payload_tval;
  wire                LsuL1_lockPort_valid;
  wire       [31:0]   LsuL1_lockPort_address;
  reg                 LsuL1_ackUnlock;
  wire                LsuL1Plugin_logic_bus_read_cmd_valid;
  wire                LsuL1Plugin_logic_bus_read_cmd_ready;
  wire       [0:0]    LsuL1Plugin_logic_bus_read_cmd_payload_id;
  wire       [31:0]   LsuL1Plugin_logic_bus_read_cmd_payload_address;
  wire                LsuL1Plugin_logic_bus_read_rsp_valid;
  wire                LsuL1Plugin_logic_bus_read_rsp_ready;
  wire       [0:0]    LsuL1Plugin_logic_bus_read_rsp_payload_id;
  wire       [255:0]  LsuL1Plugin_logic_bus_read_rsp_payload_data;
  wire                LsuL1Plugin_logic_bus_read_rsp_payload_error;
  wire                LsuL1Plugin_logic_bus_write_cmd_valid;
  wire                LsuL1Plugin_logic_bus_write_cmd_ready;
  wire                LsuL1Plugin_logic_bus_write_cmd_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  wire       [255:0]  LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  wire       [0:0]    LsuL1Plugin_logic_bus_write_cmd_payload_fragment_id;
  wire                LsuL1Plugin_logic_bus_write_rsp_valid;
  wire                LsuL1Plugin_logic_bus_write_rsp_payload_error;
  wire       [0:0]    LsuL1Plugin_logic_bus_write_rsp_payload_id;
  reg        [1:0]    LsuL1Plugin_logic_refillCompletions;
  wire                LsuL1Plugin_logic_writebackBusy;
  reg        [1:0]    LsuL1Plugin_logic_banksWrite_mask;
  reg        [6:0]    LsuL1Plugin_logic_banksWrite_address;
  reg        [255:0]  LsuL1Plugin_logic_banksWrite_writeData;
  reg        [31:0]   LsuL1Plugin_logic_banksWrite_writeMask;
  reg        [1:0]    LsuL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    LsuL1Plugin_logic_waysWrite_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_loaded;
  reg        [19:0]   LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_fault;
  wire                LsuL1Plugin_logic_waysWrite_valid;
  wire                LsuL1Plugin_logic_banks_0_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_0_write_valid;
  wire       [6:0]    LsuL1Plugin_logic_banks_0_write_payload_address;
  wire       [255:0]  LsuL1Plugin_logic_banks_0_write_payload_data;
  wire       [31:0]   LsuL1Plugin_logic_banks_0_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_0_read_cmd_valid;
  reg        [6:0]    LsuL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [255:0]  LsuL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_1_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_1_write_valid;
  wire       [6:0]    LsuL1Plugin_logic_banks_1_write_payload_address;
  wire       [255:0]  LsuL1Plugin_logic_banks_1_write_payload_data;
  wire       [31:0]   LsuL1Plugin_logic_banks_1_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_1_read_cmd_valid;
  reg        [6:0]    LsuL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [255:0]  LsuL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_0_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_1_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  reg                 LsuL1Plugin_logic_shared_write_valid;
  reg        [5:0]    LsuL1Plugin_logic_shared_write_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg        [1:0]    LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire                LsuL1Plugin_logic_shared_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_shared_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_dirty /* synthesis syn_keep = 1 */ ;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
  reg                 LsuL1Plugin_logic_refill_slots_0_valid;
  reg                 LsuL1Plugin_logic_refill_slots_0_dirty;
  reg        [31:0]   LsuL1Plugin_logic_refill_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_way;
  reg                 LsuL1Plugin_logic_refill_slots_0_cmdSent;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_priority;
  reg                 LsuL1Plugin_logic_refill_slots_0_loadedSet;
  reg                 LsuL1Plugin_logic_refill_slots_0_loaded;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_loadedCounter;
  wire                LsuL1Plugin_logic_refill_slots_0_loadedDone;
  wire                LsuL1Plugin_logic_refill_slots_0_free;
  wire                LsuL1Plugin_logic_refill_slots_0_fire;
  reg        [1:0]    LsuL1Plugin_logic_refill_slots_0_victim;
  reg                 LsuL1Plugin_logic_refill_slots_1_valid;
  reg                 LsuL1Plugin_logic_refill_slots_1_dirty;
  reg        [31:0]   LsuL1Plugin_logic_refill_slots_1_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_1_way;
  reg                 LsuL1Plugin_logic_refill_slots_1_cmdSent;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_1_priority;
  reg                 LsuL1Plugin_logic_refill_slots_1_loadedSet;
  reg                 LsuL1Plugin_logic_refill_slots_1_loaded;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_1_loadedCounter;
  wire                LsuL1Plugin_logic_refill_slots_1_loadedDone;
  wire                LsuL1Plugin_logic_refill_slots_1_free;
  wire                LsuL1Plugin_logic_refill_slots_1_fire;
  reg        [1:0]    LsuL1Plugin_logic_refill_slots_1_victim;
  wire       [1:0]    _zz_LsuL1Plugin_logic_refill_free;
  wire       [1:0]    LsuL1Plugin_logic_refill_free;
  wire                LsuL1Plugin_logic_refill_full;
  reg                 LsuL1Plugin_logic_refill_push_valid;
  wire       [31:0]   LsuL1Plugin_logic_refill_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_way;
  reg        [1:0]    LsuL1Plugin_logic_refill_push_payload_victim;
  wire                LsuL1Plugin_logic_refill_push_payload_dirty;
  wire                LsuL1Plugin_logic_refill_push_payload_unique;
  wire                LsuL1Plugin_logic_refill_push_payload_data;
  reg        [31:0]   LsuL1Plugin_logic_refill_pushCounter;
  wire                when_LsuL1Plugin_l377;
  wire                when_LsuL1Plugin_l381;
  wire                when_LsuL1Plugin_l377_1;
  wire                when_LsuL1Plugin_l381_1;
  wire                LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  wire                LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    LsuL1Plugin_logic_refill_read_arbiter_hits;
  wire                LsuL1Plugin_logic_refill_read_arbiter_hit;
  reg        [1:0]    LsuL1Plugin_logic_refill_read_arbiter_oh;
  wire                _zz_LsuL1Plugin_logic_refill_read_arbiter_sel;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_arbiter_sel;
  reg        [1:0]    LsuL1Plugin_logic_refill_read_arbiter_lock;
  wire                when_LsuL1Plugin_l301;
  wire                LsuL1Plugin_logic_bus_read_cmd_fire;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_cmdAddress;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_rspAddress;
  wire                LsuL1Plugin_logic_refill_read_dirty;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_way;
  (* keep , syn_keep *) reg        [0:0]    LsuL1Plugin_logic_refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_refill_read_rspWithData;
  reg        [1:0]    LsuL1Plugin_logic_refill_read_bankWriteNotif;
  wire                LsuL1Plugin_logic_refill_read_writeReservation_win;
  reg                 LsuL1Plugin_logic_refill_read_writeReservation_take;
  reg                 LsuL1Plugin_logic_refill_read_hadError;
  wire                when_LsuL1Plugin_l450;
  reg                 LsuL1Plugin_logic_refill_read_fire;
  wire                LsuL1Plugin_logic_refill_read_reservation_win;
  reg                 LsuL1Plugin_logic_refill_read_reservation_take;
  wire                LsuL1Plugin_logic_refill_read_faulty;
  wire                when_LsuL1Plugin_l463;
  wire       [1:0]    LsuL1_REFILL_BUSY;
  reg                 LsuL1Plugin_logic_writeback_slots_0_fire;
  reg                 LsuL1Plugin_logic_writeback_slots_0_valid;
  reg                 LsuL1Plugin_logic_writeback_slots_0_busy;
  reg        [31:0]   LsuL1Plugin_logic_writeback_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_way;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_priority;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readCmdDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readRspDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_victimBufferReady;
  reg                 LsuL1Plugin_logic_writeback_slots_0_writeCmdDone;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_timer_counter;
  wire                LsuL1Plugin_logic_writeback_slots_0_timer_done;
  wire                when_LsuL1Plugin_l530;
  wire                LsuL1Plugin_logic_writeback_slots_0_free;
  reg                 LsuL1Plugin_logic_writeback_slots_1_fire;
  reg                 LsuL1Plugin_logic_writeback_slots_1_valid;
  reg                 LsuL1Plugin_logic_writeback_slots_1_busy;
  reg        [31:0]   LsuL1Plugin_logic_writeback_slots_1_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_1_way;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_1_priority;
  reg                 LsuL1Plugin_logic_writeback_slots_1_readCmdDone;
  reg                 LsuL1Plugin_logic_writeback_slots_1_readRspDone;
  reg                 LsuL1Plugin_logic_writeback_slots_1_victimBufferReady;
  reg                 LsuL1Plugin_logic_writeback_slots_1_writeCmdDone;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_1_timer_counter;
  wire                LsuL1Plugin_logic_writeback_slots_1_timer_done;
  wire                when_LsuL1Plugin_l530_1;
  wire                LsuL1Plugin_logic_writeback_slots_1_free;
  wire       [1:0]    LsuL1_WRITEBACK_BUSY;
  wire       [1:0]    _zz_LsuL1Plugin_logic_writeback_free;
  wire       [1:0]    LsuL1Plugin_logic_writeback_free;
  wire                LsuL1Plugin_logic_writeback_full;
  reg                 LsuL1Plugin_logic_writeback_push_valid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_push_payload_way;
  wire                when_LsuL1Plugin_l556;
  wire                when_LsuL1Plugin_l561;
  wire                when_LsuL1Plugin_l556_1;
  wire                when_LsuL1Plugin_l561_1;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    LsuL1Plugin_logic_writeback_read_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_hit;
  reg        [1:0]    LsuL1Plugin_logic_writeback_read_arbiter_oh;
  wire                _zz_LsuL1Plugin_logic_writeback_read_arbiter_sel;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_sel;
  reg        [1:0]    LsuL1Plugin_logic_writeback_read_arbiter_lock;
  wire                when_LsuL1Plugin_l301_1;
  wire       [31:0]   LsuL1Plugin_logic_writeback_read_address;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_way;
  (* keep , syn_keep *) reg        [0:0]    LsuL1Plugin_logic_writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_valid;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_id;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
  wire                when_LsuL1Plugin_l605;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_valid;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_id;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way;
  wire       [255:0]  LsuL1Plugin_logic_writeback_read_readedData;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_1_0;
  wire       [1:0]    LsuL1Plugin_logic_writeback_write_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_hit;
  reg        [1:0]    LsuL1Plugin_logic_writeback_write_arbiter_oh;
  wire                _zz_LsuL1Plugin_logic_writeback_write_arbiter_sel;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_sel;
  reg        [1:0]    LsuL1Plugin_logic_writeback_write_arbiter_lock;
  wire                when_LsuL1Plugin_l301_2;
  (* keep , syn_keep *) reg        [0:0]    LsuL1Plugin_logic_writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_write_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_valid;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_ready;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_bufferRead_payload_id;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_fire;
  wire                when_LsuL1Plugin_l676;
  wire                LsuL1Plugin_logic_writeback_write_cmd_valid;
  wire                LsuL1Plugin_logic_writeback_write_cmd_ready;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_cmd_payload_id;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_bufferRead_rData_id;
  reg        [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  wire                when_Stream_l477;
  wire       [1:0]    _zz_LsuL1Plugin_logic_writeback_write_word;
  wire       [255:0]  LsuL1Plugin_logic_writeback_write_word;
  wire       [6:0]    LsuL1Plugin_logic_lsu_rb0_readAddress;
  wire                when_LsuL1Plugin_l718;
  wire                when_LsuL1Plugin_l719;
  wire                when_LsuL1Plugin_l718_1;
  wire                when_LsuL1Plugin_l719_1;
  wire                execute_lane0_ctrls_3_upIsCancel;
  wire                execute_lane0_ctrls_3_downIsCancel;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg;
  wire                when_LsuL1Plugin_l735;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg;
  wire                when_LsuL1Plugin_l735_1;
  wire                execute_lane0_ctrls_4_upIsCancel;
  wire                execute_lane0_ctrls_4_downIsCancel;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  wire                LsuL1Plugin_logic_lsu_sharedBypassers_0_hit;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  reg        [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state;
  wire                LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win;
  reg                 LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_refillHazards;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_writebackHazards;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_writebackHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_wasDirty;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty;
  wire                LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankNotRead;
  wire                LsuL1Plugin_logic_lsu_ctrl_loadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_storeHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_preventSideEffects;
  wire                LsuL1Plugin_logic_lsu_ctrl_flushHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_coherencyHazard;
  reg                 LsuL1Plugin_logic_lsu_ctrl_hazardReg;
  reg                 LsuL1Plugin_logic_lsu_ctrl_flushHazardReg;
  wire                LsuL1Plugin_logic_lsu_ctrl_canRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_canFlush;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  wire       [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1;
  reg        [1:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire                LsuL1Plugin_logic_lsu_ctrl_isAccess;
  wire                LsuL1Plugin_logic_lsu_ctrl_askRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_askUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_askFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_askCbm;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_doUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_doFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_doWrite;
  wire                LsuL1Plugin_logic_lsu_ctrl_doCbm;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_wayId;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_targetWay;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
  wire                when_LsuL1Plugin_l915;
  wire       [2:0]    _zz_23;
  wire       [3:0]    _zz_24;
  wire                when_LsuL1Plugin_l929;
  wire                when_LsuL1Plugin_l929_1;
  wire       [19:0]   _zz_LsuL1Plugin_logic_waysWrite_tag_address;
  wire                when_LsuL1Plugin_l1018;
  wire                when_LsuL1Plugin_l1025;
  wire                when_LsuL1Plugin_l1029;
  wire                when_LsuL1Plugin_l1029_1;
  wire                when_LsuL1Plugin_l1029_2;
  wire                when_LsuL1Plugin_l1029_3;
  wire                when_LsuL1Plugin_l1029_4;
  wire                when_LsuL1Plugin_l1029_5;
  wire                when_LsuL1Plugin_l1029_6;
  wire                when_LsuL1Plugin_l1029_7;
  wire                when_LsuL1Plugin_l1025_1;
  wire                when_LsuL1Plugin_l1029_8;
  wire                when_LsuL1Plugin_l1029_9;
  wire                when_LsuL1Plugin_l1029_10;
  wire                when_LsuL1Plugin_l1029_11;
  wire                when_LsuL1Plugin_l1029_12;
  wire                when_LsuL1Plugin_l1029_13;
  wire                when_LsuL1Plugin_l1029_14;
  wire                when_LsuL1Plugin_l1029_15;
  reg        [6:0]    LsuL1Plugin_logic_initializer_counter;
  wire                LsuL1Plugin_logic_initializer_done;
  wire                when_LsuL1Plugin_l1218;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg                 PrefetcherRptPlugin_logic_csr_disable;
  reg                 PrefetcherRptPlugin_logic_order_valid;
  wire                PrefetcherRptPlugin_logic_order_ready;
  wire       [31:0]   PrefetcherRptPlugin_logic_order_payload_address;
  wire                PrefetcherRptPlugin_logic_order_payload_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_payload_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_order_payload_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_order_payload_stride;
  wire                PrefetcherRptPlugin_logic_queued_valid;
  wire                PrefetcherRptPlugin_logic_queued_ready;
  wire       [31:0]   PrefetcherRptPlugin_logic_queued_payload_address;
  wire                PrefetcherRptPlugin_logic_queued_payload_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_queued_payload_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_queued_payload_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_queued_payload_stride;
  reg        [2:0]    PrefetcherRptPlugin_logic_counter;
  wire       [2:0]    PrefetcherRptPlugin_logic_advanceAt;
  wire                PrefetcherRptPlugin_logic_done;
  wire                PrefetcherRptPlugin_logic_queued_forkSerial_next_valid;
  wire                PrefetcherRptPlugin_logic_queued_forkSerial_next_ready;
  wire       [31:0]   PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_address;
  wire                PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_stride;
  wire                PrefetcherRptPlugin_logic_pip2_result_serialized_valid;
  wire                PrefetcherRptPlugin_logic_pip2_result_serialized_ready;
  wire       [31:0]   PrefetcherRptPlugin_logic_pip2_result_serialized_payload_address;
  wire                PrefetcherRptPlugin_logic_pip2_result_serialized_payload_unique;
  wire                when_StageLink_l71;
  reg                 _zz_25;
  wire                PrefetcherRptPlugin_logic_storage_read_cmd_valid;
  wire       [6:0]    PrefetcherRptPlugin_logic_storage_read_cmd_payload;
  wire       [14:0]   PrefetcherRptPlugin_logic_storage_read_rsp_tag;
  wire       [15:0]   PrefetcherRptPlugin_logic_storage_read_rsp_address;
  wire       [11:0]   PrefetcherRptPlugin_logic_storage_read_rsp_stride;
  wire       [4:0]    PrefetcherRptPlugin_logic_storage_read_rsp_score;
  wire       [2:0]    PrefetcherRptPlugin_logic_storage_read_rsp_advance;
  wire                PrefetcherRptPlugin_logic_storage_read_rsp_missed;
  wire       [51:0]   _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag;
  reg                 PrefetcherRptPlugin_logic_storage_write_valid;
  wire       [6:0]    PrefetcherRptPlugin_logic_storage_write_payload_address;
  reg        [14:0]   PrefetcherRptPlugin_logic_storage_write_payload_data_tag;
  wire       [15:0]   PrefetcherRptPlugin_logic_storage_write_payload_data_address;
  reg        [11:0]   PrefetcherRptPlugin_logic_storage_write_payload_data_stride;
  reg        [4:0]    PrefetcherRptPlugin_logic_storage_write_payload_data_score;
  reg        [2:0]    PrefetcherRptPlugin_logic_storage_write_payload_data_advance;
  wire                PrefetcherRptPlugin_logic_storage_write_payload_data_missed;
  wire                early0_MulPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_MulPlugin_logic_formatBus_payload;
  wire                early0_DivPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_DivPlugin_logic_formatBus_payload;
  wire                CsrAccessPlugin_logic_wbWi_valid;
  wire       [31:0]   CsrAccessPlugin_logic_wbWi_payload;
  reg                 CsrAccessPlugin_logic_flushPort_valid;
  reg                 PrivilegedPlugin_logic_harts_0_xretAwayFromMachine;
  wire       [1:0]    PrivilegedPlugin_logic_harts_0_commitMask;
  reg                 PrivilegedPlugin_logic_harts_0_int_pending;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_privilege;
  wire                PrivilegedPlugin_logic_harts_0_withMachinePrivilege;
  wire                PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege;
  wire                PrivilegedPlugin_logic_harts_0_hartRunning;
  wire                PrivilegedPlugin_logic_harts_0_debugMode;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mie;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mpie;
  wire       [1:0]    PrivilegedPlugin_logic_harts_0_m_status_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_fs;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_sd;
  wire                PrivilegedPlugin_logic_harts_0_m_status_tw;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mprv;
  wire                when_PrivilegedPlugin_l549;
  wire                when_PrivilegedPlugin_l550;
  wire                when_PrivilegedPlugin_l554;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  reg                 PrivilegedPlugin_logic_harts_0_m_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_m_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_meip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_mtip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_msip;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_meie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_mtie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_msie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  wire                _zz_when_TrapPlugin_l207;
  wire                _zz_when_TrapPlugin_l207_1;
  wire                _zz_when_TrapPlugin_l207_2;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready;
  reg                 TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid;
  wire                TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready;
  reg                 early0_EnvPlugin_logic_trapPort_valid;
  reg                 early0_EnvPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   early0_EnvPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    early0_EnvPlugin_logic_trapPort_payload_code;
  reg        [1:0]    early0_EnvPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    early0_EnvPlugin_logic_trapPort_payload_laneAge;
  reg                 early0_EnvPlugin_logic_flushPort_valid;
  wire                late0_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   late0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   late0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   late0_IntAluPlugin_logic_alu_result;
  wire                late0_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    late0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_patched;
  wire                late0_BranchPlugin_logic_wb_valid;
  wire       [31:0]   late0_BranchPlugin_logic_wb_payload;
  wire                late0_BranchPlugin_logic_pcPort_valid;
  wire                late0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   late0_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    late0_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid;
  wire                late0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   late0_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    late0_BranchPlugin_logic_historyPort_payload_age;
  wire                late0_BranchPlugin_logic_flushPort_valid;
  wire       [0:0]    execute_lane1_logic_trapPending;
  wire                early1_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   early1_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   early1_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   early1_IntAluPlugin_logic_alu_result;
  wire                early1_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    early1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_patched;
  wire                early1_BranchPlugin_logic_wb_valid;
  wire       [31:0]   early1_BranchPlugin_logic_wb_payload;
  wire                early1_BranchPlugin_logic_pcPort_valid;
  wire                early1_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   early1_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    early1_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid;
  wire                early1_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early1_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    early1_BranchPlugin_logic_historyPort_payload_age;
  wire                early1_BranchPlugin_logic_flushPort_valid;
  wire                late1_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   late1_IntAluPlugin_logic_wb_payload;
  wire                execute_lane1_ctrls_4_upIsCancel;
  wire                execute_lane1_ctrls_4_downIsCancel;
  (* keep , syn_keep *) reg        [31:0]   late1_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   late1_IntAluPlugin_logic_alu_result;
  wire                late1_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    late1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_patched;
  wire                late1_BranchPlugin_logic_wb_valid;
  wire       [31:0]   late1_BranchPlugin_logic_wb_payload;
  wire                late1_BranchPlugin_logic_pcPort_valid;
  wire                late1_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   late1_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    late1_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid;
  wire                late1_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   late1_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    late1_BranchPlugin_logic_historyPort_payload_age;
  wire                late1_BranchPlugin_logic_flushPort_valid;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  wire       [0:0]    FpuUnpackerPlugin_logic_packPort_cmd_at;
  reg        [1:0]    FpuUnpackerPlugin_logic_packPort_cmd_value_mode;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_value_sign;
  wire       [5:0]    FpuUnpackerPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuUnpackerPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuUnpackerPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuUnpackerPlugin_logic_packPort_cmd_roundMode;
  wire       [0:0]    FpuAddPlugin_logic_addPort_cmd_at;
  wire       [1:0]    FpuAddPlugin_logic_addPort_cmd_rs1_mode;
  wire                FpuAddPlugin_logic_addPort_cmd_rs1_quiet;
  wire                FpuAddPlugin_logic_addPort_cmd_rs1_sign;
  wire       [11:0]   FpuAddPlugin_logic_addPort_cmd_rs1_exponent;
  wire       [51:0]   FpuAddPlugin_logic_addPort_cmd_rs1_mantissa;
  wire       [1:0]    FpuAddPlugin_logic_addPort_cmd_rs2_mode;
  wire                FpuAddPlugin_logic_addPort_cmd_rs2_quiet;
  wire                FpuAddPlugin_logic_addPort_cmd_rs2_sign;
  wire       [11:0]   FpuAddPlugin_logic_addPort_cmd_rs2_exponent;
  wire       [51:0]   FpuAddPlugin_logic_addPort_cmd_rs2_mantissa;
  wire       [0:0]    FpuAddPlugin_logic_addPort_cmd_format;
  wire       [2:0]    FpuAddPlugin_logic_addPort_cmd_roundMode;
  wire       [0:0]    FpuMulPlugin_logic_packPort_cmd_at;
  wire       [1:0]    FpuMulPlugin_logic_packPort_cmd_value_mode;
  wire                FpuMulPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuMulPlugin_logic_packPort_cmd_value_sign;
  wire       [12:0]   FpuMulPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuMulPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuMulPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuMulPlugin_logic_packPort_cmd_roundMode;
  wire       [0:0]    FpuSqrtPlugin_logic_packPort_cmd_at;
  reg        [1:0]    FpuSqrtPlugin_logic_packPort_cmd_value_mode;
  reg                 FpuSqrtPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuSqrtPlugin_logic_packPort_cmd_value_sign;
  wire       [10:0]   FpuSqrtPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuSqrtPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuSqrtPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuSqrtPlugin_logic_packPort_cmd_roundMode;
  wire                FpuClassPlugin_logic_iwb_valid;
  wire       [31:0]   FpuClassPlugin_logic_iwb_payload;
  wire                FpuCmpPlugin_logic_ffwb_flags_NX;
  wire                FpuCmpPlugin_logic_ffwb_flags_UF;
  wire                FpuCmpPlugin_logic_ffwb_flags_OF;
  wire                FpuCmpPlugin_logic_ffwb_flags_DZ;
  wire                FpuCmpPlugin_logic_ffwb_flags_NV;
  wire       [0:0]    FpuCmpPlugin_logic_ffwb_ats;
  wire                FpuCmpPlugin_logic_fwb_valid;
  reg        [63:0]   FpuCmpPlugin_logic_fwb_payload;
  wire                FpuCmpPlugin_logic_iwb_valid;
  wire       [31:0]   FpuCmpPlugin_logic_iwb_payload;
  wire                FpuF2iPlugin_logic_ffwb_flags_NX;
  wire                FpuF2iPlugin_logic_ffwb_flags_UF;
  wire                FpuF2iPlugin_logic_ffwb_flags_OF;
  wire                FpuF2iPlugin_logic_ffwb_flags_DZ;
  wire                FpuF2iPlugin_logic_ffwb_flags_NV;
  wire       [0:0]    FpuF2iPlugin_logic_ffwb_ats;
  wire                FpuF2iPlugin_logic_iwb_valid;
  wire       [31:0]   FpuF2iPlugin_logic_iwb_payload;
  wire                FpuMvPlugin_logic_fwb_valid;
  reg        [63:0]   FpuMvPlugin_logic_fwb_payload;
  wire                FpuMvPlugin_logic_iwb_valid;
  wire       [31:0]   FpuMvPlugin_logic_iwb_payload;
  wire       [0:0]    FpuXxPlugin_logic_packPort_cmd_at;
  wire       [1:0]    FpuXxPlugin_logic_packPort_cmd_value_mode;
  wire                FpuXxPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuXxPlugin_logic_packPort_cmd_value_sign;
  wire       [11:0]   FpuXxPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuXxPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuXxPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuXxPlugin_logic_packPort_cmd_roundMode;
  wire       [0:0]    FpuDivPlugin_logic_packPort_cmd_at;
  reg        [1:0]    FpuDivPlugin_logic_packPort_cmd_value_mode;
  reg                 FpuDivPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuDivPlugin_logic_packPort_cmd_value_sign;
  wire       [12:0]   FpuDivPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuDivPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuDivPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuDivPlugin_logic_packPort_cmd_roundMode;
  wire                WhiteboxerPlugin_logic_fetch_fire;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_valid;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_last;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_write;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_id;
  wire       [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_address;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_valid;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_last;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_write;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_id;
  wire       [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_address;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_valid;
  reg                 LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_last;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_write;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_id;
  reg        [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_address;
  wire       [255:0]  LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_data;
  reg        [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_counter;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_fire;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_ready;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_last;
  wire                LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_write;
  wire       [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_id;
  wire       [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_address;
  wire       [255:0]  LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_data;
  reg                 LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rValid;
  reg                 LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_last;
  reg                 LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_write;
  reg        [0:0]    LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_id;
  reg        [31:0]   LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_address;
  reg        [255:0]  LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_data;
  wire                when_Stream_l477_1;
  reg        [3:0]    CsrAccessPlugin_bus_decode_trapCode;
  wire                CsrAccessPlugin_bus_read_valid;
  wire                CsrAccessPlugin_bus_read_moving;
  wire       [11:0]   CsrAccessPlugin_bus_read_address;
  reg                 CsrAccessPlugin_bus_read_halt;
  wire       [31:0]   CsrAccessPlugin_bus_read_toWriteBits;
  wire       [31:0]   CsrAccessPlugin_bus_read_data;
  wire                CsrAccessPlugin_bus_write_valid;
  wire                CsrAccessPlugin_bus_write_moving;
  reg                 CsrAccessPlugin_bus_write_halt;
  reg        [31:0]   CsrAccessPlugin_bus_write_bits;
  wire       [11:0]   CsrAccessPlugin_bus_write_address;
  reg        [3:0]    FetchL1Plugin_logic_trapPort_payload_code;
  reg        [1:0]    FetchL1Plugin_logic_trapPort_payload_arg;
  wire                FetchL1Plugin_logic_banks_0_write_valid;
  wire       [6:0]    FetchL1Plugin_logic_banks_0_write_payload_address;
  wire       [255:0]  FetchL1Plugin_logic_banks_0_write_payload_data;
  wire                FetchL1Plugin_logic_banks_0_read_cmd_valid;
  wire       [6:0]    FetchL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [255:0]  FetchL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_banks_1_write_valid;
  wire       [6:0]    FetchL1Plugin_logic_banks_1_write_payload_address;
  wire       [255:0]  FetchL1Plugin_logic_banks_1_write_payload_data;
  wire                FetchL1Plugin_logic_banks_1_read_cmd_valid;
  wire       [6:0]    FetchL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [255:0]  FetchL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [1:0]    FetchL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    FetchL1Plugin_logic_waysWrite_address;
  reg                 FetchL1Plugin_logic_waysWrite_tag_loaded;
  reg                 FetchL1Plugin_logic_waysWrite_tag_error;
  reg        [19:0]   FetchL1Plugin_logic_waysWrite_tag_address;
  wire                FetchL1Plugin_logic_ways_0_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_1_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_1_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_1_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  reg                 FetchL1Plugin_logic_plru_write_valid;
  reg        [5:0]    FetchL1Plugin_logic_plru_write_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_plru_write_payload_data_0;
  wire                FetchL1Plugin_logic_plru_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_plru_read_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    FetchL1Plugin_logic_plru_read_rsp_0 /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_invalidate_cmd_valid;
  wire                FetchL1Plugin_logic_invalidate_cmd_ready;
  reg                 FetchL1Plugin_logic_invalidate_canStart;
  reg        [6:0]    FetchL1Plugin_logic_invalidate_counter;
  wire       [6:0]    FetchL1Plugin_logic_invalidate_counterIncr;
  wire                FetchL1Plugin_logic_invalidate_done;
  wire                FetchL1Plugin_logic_invalidate_last;
  reg                 FetchL1Plugin_logic_invalidate_firstEver;
  wire                when_FetchL1Plugin_l204;
  wire                when_FetchL1Plugin_l211;
  wire                when_FetchL1Plugin_l216;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  reg                 FetchL1Plugin_logic_refill_start_valid;
  wire       [31:0]   FetchL1Plugin_logic_refill_start_address;
  wire       [0:0]    FetchL1Plugin_logic_refill_start_wayToAllocate;
  wire                FetchL1Plugin_logic_refill_start_isIo;
  reg                 FetchL1Plugin_logic_refill_slots_0_valid;
  reg                 FetchL1Plugin_logic_refill_slots_0_cmdSent;
  (* keep , syn_keep *) reg        [31:0]   FetchL1Plugin_logic_refill_slots_0_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_refill_slots_0_isIo;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  reg        [1:0]    FetchL1Plugin_logic_refill_slots_0_priority;
  wire                FetchL1Plugin_logic_refill_slots_0_askCmd;
  reg                 FetchL1Plugin_logic_refill_slots_1_valid;
  reg                 FetchL1Plugin_logic_refill_slots_1_cmdSent;
  (* keep , syn_keep *) reg        [31:0]   FetchL1Plugin_logic_refill_slots_1_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_refill_slots_1_isIo;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_1_wayToAllocate;
  reg        [1:0]    FetchL1Plugin_logic_refill_slots_1_priority;
  wire                FetchL1Plugin_logic_refill_slots_1_askCmd;
  wire                when_FetchL1Plugin_l246;
  wire                when_FetchL1Plugin_l246_1;
  reg        [31:0]   FetchL1Plugin_logic_refill_pushCounter;
  wire                _zz_38;
  wire       [1:0]    _zz_39;
  wire                FetchL1Plugin_logic_refill_hazard;
  wire                when_FetchL1Plugin_l255;
  wire                when_FetchL1Plugin_l268;
  wire       [1:0]    FetchL1Plugin_logic_refill_onCmd_propoedOh;
  reg                 FetchL1Plugin_logic_refill_onCmd_locked;
  wire                when_FetchL1Plugin_l276;
  reg        [1:0]    FetchL1Plugin_logic_refill_onCmd_lockedOh;
  wire       [1:0]    FetchL1Plugin_logic_refill_onCmd_oh;
  wire                _zz_FetchL1Plugin_logic_bus_cmd_payload_address;
  wire                _zz_FetchL1Plugin_logic_bus_cmd_payload_id;
  reg        [0:0]    FetchL1Plugin_logic_refill_onRsp_rspIdReg;
  (* keep , syn_keep *) reg        [0:0]    FetchL1Plugin_logic_refill_onRsp_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_refill_onRsp_holdHarts;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297;
  reg                 FetchL1Plugin_logic_refill_onRsp_firstCycle;
  wire                FetchL1Plugin_logic_bus_rsp_fire;
  wire       [0:0]    FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  wire       [31:0]   FetchL1Plugin_logic_refill_onRsp_address;
  wire                when_FetchL1Plugin_l304;
  wire                when_FetchL1Plugin_l330;
  wire                FetchL1Plugin_logic_cmd_doIt;
  wire       [31:0]   FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
  wire       [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
  reg                 FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
  reg        [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
  wire                FetchL1Plugin_logic_ctrl_dataAccessFault;
  reg                 FetchL1Plugin_logic_ctrl_trapSent;
  reg                 FetchL1Plugin_logic_ctrl_allowRefill;
  wire                when_FetchL1Plugin_l474;
  wire                when_FetchL1Plugin_l480;
  wire                when_FetchL1Plugin_l487;
  wire                when_FetchL1Plugin_l520;
  wire                when_FetchL1Plugin_l533;
  wire                when_FetchL1Plugin_l537;
  reg                 FetchL1Plugin_logic_ctrl_firstCycle;
  wire                when_FetchL1Plugin_l541;
  wire                when_FetchL1Plugin_l558;
  reg        [3:0]    LsuPlugin_logic_trapPort_payload_code;
  reg        [1:0]    LsuPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    LsuPlugin_logic_trapPort_payload_laneAge;
  reg                 LsuPlugin_logic_flushPort_valid;
  wire       [15:0]   LsuPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    LsuPlugin_logic_flushPort_payload_laneAge;
  wire                LsuPlugin_logic_flushPort_payload_self;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_0;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_1;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_2;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_3;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_4;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_5;
  wire                LsuPlugin_logic_commitProbe_valid;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_pc;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_address;
  wire                LsuPlugin_logic_commitProbe_payload_load;
  wire                LsuPlugin_logic_commitProbe_payload_store;
  wire                LsuPlugin_logic_commitProbe_payload_trap;
  wire                LsuPlugin_logic_commitProbe_payload_io;
  wire                LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  wire                LsuPlugin_logic_commitProbe_payload_miss;
  wire                LsuPlugin_logic_iwb_valid;
  reg        [31:0]   LsuPlugin_logic_iwb_payload;
  wire                execute_lane0_ctrls_0_upIsCancel;
  wire                execute_lane0_ctrls_0_downIsCancel;
  wire                GSharePlugin_logic_mem_write_valid;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_1;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_2;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_3;
  wire                GSharePlugin_logic_mem_writes_0_valid;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_0;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_1;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_2;
  wire       [1:0]    GSharePlugin_logic_mem_writes_0_payload_data_3;
  wire       [1:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  wire       [1:0]    _zz_GSharePlugin_logic_readRsp_readed_0_0;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_0;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_1;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_2;
  wire       [1:0]    GSharePlugin_logic_readRsp_readed_0_3;
  wire       [7:0]    _zz_GSharePlugin_logic_readRsp_readed_0_0_1;
  wire                when_GSharePlugin_l100;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_push;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop;
  reg                 BtbPlugin_logic_ras_ptr_pushIt;
  reg                 BtbPlugin_logic_ras_ptr_popIt;
  wire                BtbPlugin_logic_ras_readIt;
  reg        [30:0]   BtbPlugin_logic_ras_read;
  wire                BtbPlugin_logic_ras_write_valid;
  wire       [1:0]    BtbPlugin_logic_ras_write_payload_address;
  reg        [30:0]   BtbPlugin_logic_ras_write_payload_data;
  reg                 BtbPlugin_logic_memWrite_valid;
  reg        [6:0]    BtbPlugin_logic_memWrite_payload_address;
  reg        [11:0]   BtbPlugin_logic_memWrite_payload_data_0_hash;
  reg        [0:0]    BtbPlugin_logic_memWrite_payload_data_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPush;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPop;
  reg        [11:0]   BtbPlugin_logic_memWrite_payload_data_1_hash;
  reg        [0:0]    BtbPlugin_logic_memWrite_payload_data_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memWrite_payload_data_1_pcTarget;
  reg                 BtbPlugin_logic_memWrite_payload_data_1_isBranch;
  reg                 BtbPlugin_logic_memWrite_payload_data_1_isPush;
  reg                 BtbPlugin_logic_memWrite_payload_data_1_isPop;
  reg        [1:0]    BtbPlugin_logic_memWrite_payload_mask;
  wire                BtbPlugin_logic_memRead_cmd_valid;
  wire       [6:0]    BtbPlugin_logic_memRead_cmd_payload;
  wire       [11:0]   BtbPlugin_logic_memRead_rsp_0_hash;
  wire       [0:0]    BtbPlugin_logic_memRead_rsp_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memRead_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memRead_rsp_0_isBranch;
  wire                BtbPlugin_logic_memRead_rsp_0_isPush;
  wire                BtbPlugin_logic_memRead_rsp_0_isPop;
  wire       [11:0]   BtbPlugin_logic_memRead_rsp_1_hash;
  wire       [0:0]    BtbPlugin_logic_memRead_rsp_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memRead_rsp_1_pcTarget;
  wire                BtbPlugin_logic_memRead_rsp_1_isBranch;
  wire                BtbPlugin_logic_memRead_rsp_1_isPush;
  wire                BtbPlugin_logic_memRead_rsp_1_isPop;
  wire                BtbPlugin_logic_memDp_wp_valid;
  wire       [6:0]    BtbPlugin_logic_memDp_wp_payload_address;
  wire       [11:0]   BtbPlugin_logic_memDp_wp_payload_data_0_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isBranch;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPush;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPop;
  wire       [11:0]   BtbPlugin_logic_memDp_wp_payload_data_1_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_wp_payload_data_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memDp_wp_payload_data_1_pcTarget;
  wire                BtbPlugin_logic_memDp_wp_payload_data_1_isBranch;
  wire                BtbPlugin_logic_memDp_wp_payload_data_1_isPush;
  wire                BtbPlugin_logic_memDp_wp_payload_data_1_isPop;
  wire       [1:0]    BtbPlugin_logic_memDp_wp_payload_mask;
  wire                BtbPlugin_logic_memDp_rp_cmd_valid;
  wire       [6:0]    BtbPlugin_logic_memDp_rp_cmd_payload;
  wire       [11:0]   BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_rp_rsp_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  wire       [11:0]   BtbPlugin_logic_memDp_rp_rsp_1_hash;
  wire       [0:0]    BtbPlugin_logic_memDp_rp_rsp_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_memDp_rp_rsp_1_pcTarget;
  wire                BtbPlugin_logic_memDp_rp_rsp_1_isBranch;
  wire                BtbPlugin_logic_memDp_rp_rsp_1_isPush;
  wire                BtbPlugin_logic_memDp_rp_rsp_1_isPop;
  wire       [93:0]   _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [46:0]   _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1;
  wire       [46:0]   _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash;
  wire       [9:0]    WhiteboxerPlugin_logic_fetch_fetchId;
  wire                WhiteboxerPlugin_logic_decodes_0_fire;
  reg                 decode_ctrls_0_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50;
  wire                WhiteboxerPlugin_logic_decodes_0_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_decodeId;
  wire                WhiteboxerPlugin_logic_decodes_1_fire;
  reg                 decode_ctrls_0_up_LANE_SEL_1_regNext;
  wire                when_CtrlLaneApi_l50_1;
  wire                WhiteboxerPlugin_logic_decodes_1_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_1_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_1_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_1_decodeId;
  wire       [15:0]   early0_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early0_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                early0_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   CsrAccessPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    CsrAccessPlugin_logic_flushPort_payload_laneAge;
  wire                CsrAccessPlugin_logic_flushPort_payload_self;
  reg                 CsrAccessPlugin_logic_trapPort_valid;
  reg                 CsrAccessPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   CsrAccessPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    CsrAccessPlugin_logic_trapPort_payload_code;
  wire       [1:0]    CsrAccessPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    CsrAccessPlugin_logic_trapPort_payload_laneAge;
  wire       [15:0]   early0_EnvPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early0_EnvPlugin_logic_flushPort_payload_laneAge;
  wire                early0_EnvPlugin_logic_flushPort_payload_self;
  wire       [15:0]   late0_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    late0_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                late0_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   early1_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early1_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                early1_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   late1_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    late1_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                late1_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   FpuUnpackerPlugin_logic_packPort_cmd_uopId;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_flags_DZ;
  wire                FpuUnpackerPlugin_logic_packPort_cmd_flags_NV;
  wire       [15:0]   FpuAddPlugin_logic_addPort_cmd_uopId;
  wire                FpuAddPlugin_logic_addPort_cmd_flags_NX;
  wire                FpuAddPlugin_logic_addPort_cmd_flags_UF;
  wire                FpuAddPlugin_logic_addPort_cmd_flags_OF;
  wire                FpuAddPlugin_logic_addPort_cmd_flags_DZ;
  wire                FpuAddPlugin_logic_addPort_cmd_flags_NV;
  wire       [15:0]   FpuMulPlugin_logic_packPort_cmd_uopId;
  wire                FpuMulPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuMulPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuMulPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuMulPlugin_logic_packPort_cmd_flags_DZ;
  wire                FpuMulPlugin_logic_packPort_cmd_flags_NV;
  wire       [0:0]    FpuMulPlugin_logic_addPort_cmd_at;
  wire       [1:0]    FpuMulPlugin_logic_addPort_cmd_rs1_mode;
  wire                FpuMulPlugin_logic_addPort_cmd_rs1_quiet;
  wire                FpuMulPlugin_logic_addPort_cmd_rs1_sign;
  wire       [12:0]   FpuMulPlugin_logic_addPort_cmd_rs1_exponent;
  wire       [104:0]  FpuMulPlugin_logic_addPort_cmd_rs1_mantissa;
  wire       [1:0]    FpuMulPlugin_logic_addPort_cmd_rs2_mode;
  wire                FpuMulPlugin_logic_addPort_cmd_rs2_quiet;
  wire                FpuMulPlugin_logic_addPort_cmd_rs2_sign;
  wire       [11:0]   FpuMulPlugin_logic_addPort_cmd_rs2_exponent;
  wire       [51:0]   FpuMulPlugin_logic_addPort_cmd_rs2_mantissa;
  wire       [0:0]    FpuMulPlugin_logic_addPort_cmd_format;
  wire       [2:0]    FpuMulPlugin_logic_addPort_cmd_roundMode;
  wire       [15:0]   FpuMulPlugin_logic_addPort_cmd_uopId;
  wire                FpuMulPlugin_logic_addPort_cmd_flags_NX;
  wire                FpuMulPlugin_logic_addPort_cmd_flags_UF;
  wire                FpuMulPlugin_logic_addPort_cmd_flags_OF;
  wire                FpuMulPlugin_logic_addPort_cmd_flags_DZ;
  wire                FpuMulPlugin_logic_addPort_cmd_flags_NV;
  wire       [15:0]   FpuSqrtPlugin_logic_packPort_cmd_uopId;
  wire                FpuSqrtPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuSqrtPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuSqrtPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuSqrtPlugin_logic_packPort_cmd_flags_DZ;
  wire                FpuSqrtPlugin_logic_packPort_cmd_flags_NV;
  wire       [15:0]   FpuXxPlugin_logic_packPort_cmd_uopId;
  wire                FpuXxPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuXxPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuXxPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuXxPlugin_logic_packPort_cmd_flags_DZ;
  wire                FpuXxPlugin_logic_packPort_cmd_flags_NV;
  wire       [15:0]   FpuDivPlugin_logic_packPort_cmd_uopId;
  wire                FpuDivPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuDivPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuDivPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuDivPlugin_logic_packPort_cmd_flags_DZ;
  reg                 FpuDivPlugin_logic_packPort_cmd_flags_NV;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l701;
  wire       [31:0]   FetchL1Plugin_pmaBuilder_addressBits;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_hit;
  wire                _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  reg        [0:0]    FetchL1Plugin_logic_bus_toWishbone_counter;
  wire                FetchL1Plugin_logic_bus_toWishbone_pending;
  wire                FetchL1Plugin_logic_bus_toWishbone_lastCycle;
  wire                when_FetchL1Bus_l247;
  wire                when_FetchL1Bus_l250;
  reg                 _zz_FetchL1Plugin_logic_bus_rsp_valid;
  reg        [0:0]    FetchL1Plugin_logic_bus_cmd_payload_id_regNext;
  reg        [255:0]  FetchL1WishbonePlugin_logic_bus_DAT_MISO_regNext;
  reg                 FetchL1WishbonePlugin_logic_bus_ERR_regNext;
  reg                 DecoderPlugin_logic_forgetPort_valid;
  reg        [31:0]   DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire                execute_lane0_ctrls_1_upIsCancel;
  wire                execute_lane0_ctrls_1_downIsCancel;
  reg        [31:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  reg        [31:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   early0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  reg        [31:0]   lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [4:0]    lane0_IntFormatPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_1_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_2_wb_payload;
  wire       [4:0]    lane0_IntFormatPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_2_raw;
  reg        [31:0]   _zz_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  reg        [31:0]   _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   late0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                execute_lane1_ctrls_1_upIsCancel;
  wire                execute_lane1_ctrls_1_downIsCancel;
  reg        [31:0]   _zz_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   early1_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane1_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [1:0]    lane1_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_0_raw;
  wire                lane1_IntFormatPlugin_logic_stages_1_wb_valid;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [1:0]    lane1_IntFormatPlugin_logic_stages_1_hits;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_1_raw;
  wire                execute_lane1_ctrls_3_upIsCancel;
  wire                execute_lane1_ctrls_3_downIsCancel;
  reg        [31:0]   _zz_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   late1_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                FpuAddSharedPlugin_logic_completion_valid;
  wire       [15:0]   FpuAddSharedPlugin_logic_completion_payload_uopId;
  wire                FpuAddSharedPlugin_logic_completion_payload_trap;
  wire                FpuAddSharedPlugin_logic_completion_payload_commit;
  wire       [1:0]    FpuAddSharedPlugin_logic_packPort_cmd_at;
  wire       [1:0]    FpuAddSharedPlugin_logic_packPort_cmd_value_mode;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_value_quiet;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_value_sign;
  wire       [12:0]   FpuAddSharedPlugin_logic_packPort_cmd_value_exponent;
  wire       [53:0]   FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa;
  wire       [0:0]    FpuAddSharedPlugin_logic_packPort_cmd_format;
  wire       [2:0]    FpuAddSharedPlugin_logic_packPort_cmd_roundMode;
  wire       [15:0]   FpuAddSharedPlugin_logic_packPort_cmd_uopId;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_flags_NX;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_flags_UF;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_flags_OF;
  wire                FpuAddSharedPlugin_logic_packPort_cmd_flags_DZ;
  reg                 FpuAddSharedPlugin_logic_packPort_cmd_flags_NV;
  wire       [1:0]    FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs1_0_quiet;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs1_0_sign;
  wire       [12:0]   FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent;
  wire       [104:0]  FpuAddSharedPlugin_logic_inserter_portsRs1_0_mantissa;
  wire       [1:0]    FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs1_1_quiet;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs1_1_sign;
  wire       [12:0]   FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent;
  wire       [104:0]  FpuAddSharedPlugin_logic_inserter_portsRs1_1_mantissa;
  wire       [1:0]    FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs2_0_quiet;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs2_0_sign;
  wire       [11:0]   FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent;
  wire       [51:0]   FpuAddSharedPlugin_logic_inserter_portsRs2_0_mantissa;
  wire       [1:0]    FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs2_1_quiet;
  wire                FpuAddSharedPlugin_logic_inserter_portsRs2_1_sign;
  wire       [11:0]   FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent;
  wire       [51:0]   FpuAddSharedPlugin_logic_inserter_portsRs2_1_mantissa;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_0_valid;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode;
  wire       [121:0]  _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode;
  wire       [67:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1;
  wire       [1:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1;
  wire       [0:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT;
  wire       [0:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1;
  wire       [2:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE;
  wire       [2:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1;
  wire       [4:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX;
  wire       [12:0]   _zz_when_AFix_l1168;
  reg        [12:0]   _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs;
  wire                when_AFix_l1168;
  reg        [6:0]    _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat;
  wire                when_UInt_l119;
  wire       [107:0]  _zz_when_Utils_l1585_14;
  reg                 _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1;
  wire                when_Utils_l1585;
  wire                when_Utils_l1585_1;
  wire                when_Utils_l1585_2;
  wire                when_Utils_l1585_3;
  wire                when_Utils_l1585_4;
  wire                when_Utils_l1585_5;
  wire                when_Utils_l1585_6;
  wire                when_FpuAdd_l56;
  wire       [106:0]  _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned;
  wire       [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_31;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_32;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_35;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_36;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_39;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_40;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_43;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_44;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_47;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_48;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_51;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_52;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_55;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_56;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_59;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_60;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_63;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_64;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_67;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_68;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_71;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_72;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_75;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_76;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_79;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_80;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_83;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_84;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_87;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_88;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_91;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_92;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_95;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_96;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_99;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_100;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_103;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_104;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_106;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_107;
  reg        [107:0]  _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_112;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_114;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_119;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_121;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_127;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_129;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_135;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_137;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_143;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_145;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_150;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_152;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_156;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_157;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_1;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_2;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_3;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_4;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_5;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_6;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_7;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_8;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_9;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_11;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_12;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_13;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_14;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_15;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_16;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_18;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_19;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_20;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_22;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_26;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_27;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_28;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_29;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_30;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_31;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_33;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_34;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_35;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_37;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_41;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_42;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_43;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_45;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_49;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_57;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_58;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_59;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_60;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_61;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_62;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_64;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_65;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_66;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_68;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_72;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_73;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_74;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_76;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_80;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_88;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_89;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_90;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_92;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_96;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105;
  wire                _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106;
  wire                when_FpuAdd_l101;
  wire                when_FpuAdd_l104;
  wire                execute_lane0_ctrls_6_upIsCancel;
  wire                execute_lane0_ctrls_6_downIsCancel;
  wire                execute_lane0_ctrls_9_upIsCancel;
  wire                execute_lane0_ctrls_9_downIsCancel;
  wire       [1:0]    FpuAddSharedPlugin_logic_onPack_mask;
  wire       [107:0]  _zz_when_AFix_l852;
  reg        [53:0]   _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa;
  wire                when_AFix_l852;
  reg                 FpuUnpackerPlugin_logic_unpacker_results_0_valid;
  wire       [5:0]    FpuUnpackerPlugin_logic_unpacker_results_0_payload_shift;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_results_0_payload_data;
  reg                 FpuUnpackerPlugin_logic_unpacker_results_1_valid;
  wire       [5:0]    FpuUnpackerPlugin_logic_unpacker_results_1_payload_shift;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_results_1_payload_data;
  wire       [52:0]   _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_12;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_15;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_16;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_19;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_20;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_23;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_24;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_27;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_28;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_31;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_32;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_35;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_36;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_39;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_40;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_43;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_44;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_47;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_48;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_51;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_52;
  reg        [52:0]   _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_57;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_59;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_64;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_66;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_72;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_74;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75;
  wire       [52:0]   _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_77;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_78;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_79;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_80;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_81;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_82;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_83;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_84;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_85;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_86;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_88;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_89;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_90;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_91;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_92;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_93;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_95;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_96;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_97;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_99;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_103;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_104;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_105;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_106;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_107;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_108;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_110;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_111;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_112;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_114;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_118;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_119;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_120;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_122;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127;
  wire                _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128;
  wire       [51:0]   FpuUnpackerPlugin_logic_unpacker_logic_shifter;
  wire       [1:0]    _zz_46;
  reg                 FpuUnpackerPlugin_logic_onUnpack_firstCycle;
  wire                when_FpuUnpackerPlugin_l165;
  reg        [2:0]    FpuUnpackerPlugin_logic_onUnpack_fsmRequesters;
  reg        [2:0]    FpuUnpackerPlugin_logic_onUnpack_fsmServed;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5;
  reg        [43:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6;
  reg        [110:0]  _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  reg        [110:0]  _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1;
  reg                 early0_DivPlugin_logic_processing_divRevertResult;
  reg                 early0_DivPlugin_logic_processing_cmdSent;
  wire                io_cmd_fire;
  reg                 early0_DivPlugin_logic_processing_request;
  reg        [63:0]   early0_DivPlugin_logic_processing_a;
  reg        [63:0]   early0_DivPlugin_logic_processing_b;
  reg                 early0_DivPlugin_logic_processing_unscheduleRequest;
  wire                early0_DivPlugin_logic_processing_freeze;
  wire       [31:0]   early0_DivPlugin_logic_processing_selected;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire       [1:0]    early0_EnvPlugin_logic_exe_privilege;
  wire       [1:0]    early0_EnvPlugin_logic_exe_xretPriv;
  reg                 early0_EnvPlugin_logic_exe_commit;
  wire                early0_EnvPlugin_logic_exe_retKo;
  wire                early0_EnvPlugin_logic_exe_vmaKo;
  wire                when_EnvPlugin_l86;
  wire                when_EnvPlugin_l95;
  wire                when_EnvPlugin_l119;
  wire                when_EnvPlugin_l123;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_a;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early0_BranchPlugin_pcCalc_slices;
  reg        [31:0]   early1_BranchPlugin_pcCalc_target_a;
  reg        [31:0]   early1_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early1_BranchPlugin_pcCalc_slices;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_0;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_1;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_2;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_3;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_0;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_1;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_2;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_3;
  wire       [15:0]   AlignerPlugin_logic_slices_data_0;
  wire       [15:0]   AlignerPlugin_logic_slices_data_1;
  wire       [15:0]   AlignerPlugin_logic_slices_data_2;
  wire       [15:0]   AlignerPlugin_logic_slices_data_3;
  wire       [15:0]   AlignerPlugin_logic_slices_data_4;
  wire       [15:0]   AlignerPlugin_logic_slices_data_5;
  wire       [15:0]   AlignerPlugin_logic_slices_data_6;
  wire       [15:0]   AlignerPlugin_logic_slices_data_7;
  wire       [7:0]    AlignerPlugin_logic_slices_mask;
  wire       [7:0]    AlignerPlugin_logic_slices_last;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_0;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_1;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_2;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_3;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_4;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_5;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_6;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_7;
  reg        [7:0]    AlignerPlugin_logic_scanners_0_usageMask;
  wire                AlignerPlugin_logic_scanners_0_checker_0_required;
  wire                AlignerPlugin_logic_scanners_0_checker_0_last;
  wire                AlignerPlugin_logic_scanners_0_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_0_present;
  wire                AlignerPlugin_logic_scanners_0_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_0_checker_1_required;
  wire                AlignerPlugin_logic_scanners_0_checker_1_last;
  wire                AlignerPlugin_logic_scanners_0_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_1_present;
  wire                AlignerPlugin_logic_scanners_0_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_0_redo;
  wire                AlignerPlugin_logic_scanners_0_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_1_usageMask;
  wire                AlignerPlugin_logic_scanners_1_checker_0_required;
  wire                AlignerPlugin_logic_scanners_1_checker_0_last;
  wire                AlignerPlugin_logic_scanners_1_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_0_present;
  wire                AlignerPlugin_logic_scanners_1_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_1_checker_1_required;
  wire                AlignerPlugin_logic_scanners_1_checker_1_last;
  wire                AlignerPlugin_logic_scanners_1_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_1_present;
  wire                AlignerPlugin_logic_scanners_1_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_1_redo;
  wire                AlignerPlugin_logic_scanners_1_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_2_usageMask;
  wire                AlignerPlugin_logic_scanners_2_checker_0_required;
  wire                AlignerPlugin_logic_scanners_2_checker_0_last;
  wire                AlignerPlugin_logic_scanners_2_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_0_present;
  wire                AlignerPlugin_logic_scanners_2_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_2_checker_1_required;
  wire                AlignerPlugin_logic_scanners_2_checker_1_last;
  wire                AlignerPlugin_logic_scanners_2_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_1_present;
  wire                AlignerPlugin_logic_scanners_2_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_2_redo;
  wire                AlignerPlugin_logic_scanners_2_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_3_usageMask;
  wire                AlignerPlugin_logic_scanners_3_checker_0_required;
  wire                AlignerPlugin_logic_scanners_3_checker_0_last;
  wire                AlignerPlugin_logic_scanners_3_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_0_present;
  wire                AlignerPlugin_logic_scanners_3_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_3_checker_1_required;
  wire                AlignerPlugin_logic_scanners_3_checker_1_last;
  wire                AlignerPlugin_logic_scanners_3_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_1_present;
  wire                AlignerPlugin_logic_scanners_3_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_3_redo;
  wire                AlignerPlugin_logic_scanners_3_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_4_usageMask;
  wire                AlignerPlugin_logic_scanners_4_checker_0_required;
  wire                AlignerPlugin_logic_scanners_4_checker_0_last;
  wire                AlignerPlugin_logic_scanners_4_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_4_checker_0_present;
  wire                AlignerPlugin_logic_scanners_4_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_4_checker_1_required;
  wire                AlignerPlugin_logic_scanners_4_checker_1_last;
  wire                AlignerPlugin_logic_scanners_4_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_4_checker_1_present;
  wire                AlignerPlugin_logic_scanners_4_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_4_redo;
  wire                AlignerPlugin_logic_scanners_4_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_5_usageMask;
  wire                AlignerPlugin_logic_scanners_5_checker_0_required;
  wire                AlignerPlugin_logic_scanners_5_checker_0_last;
  wire                AlignerPlugin_logic_scanners_5_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_5_checker_0_present;
  wire                AlignerPlugin_logic_scanners_5_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_5_checker_1_required;
  wire                AlignerPlugin_logic_scanners_5_checker_1_last;
  wire                AlignerPlugin_logic_scanners_5_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_5_checker_1_present;
  wire                AlignerPlugin_logic_scanners_5_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_5_redo;
  wire                AlignerPlugin_logic_scanners_5_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_6_usageMask;
  wire                AlignerPlugin_logic_scanners_6_checker_0_required;
  wire                AlignerPlugin_logic_scanners_6_checker_0_last;
  wire                AlignerPlugin_logic_scanners_6_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_6_checker_0_present;
  wire                AlignerPlugin_logic_scanners_6_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_6_checker_1_required;
  wire                AlignerPlugin_logic_scanners_6_checker_1_last;
  wire                AlignerPlugin_logic_scanners_6_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_6_checker_1_present;
  wire                AlignerPlugin_logic_scanners_6_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_6_redo;
  wire                AlignerPlugin_logic_scanners_6_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_7_usageMask;
  wire                AlignerPlugin_logic_scanners_7_checker_0_required;
  wire                AlignerPlugin_logic_scanners_7_checker_0_last;
  wire                AlignerPlugin_logic_scanners_7_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_7_checker_0_present;
  wire                AlignerPlugin_logic_scanners_7_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_7_checker_1_required;
  wire                AlignerPlugin_logic_scanners_7_checker_1_last;
  wire                AlignerPlugin_logic_scanners_7_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_7_checker_1_present;
  wire                AlignerPlugin_logic_scanners_7_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_7_redo;
  wire                AlignerPlugin_logic_scanners_7_valid;
  wire       [7:0]    AlignerPlugin_logic_usedMask_0;
  wire       [7:0]    AlignerPlugin_logic_usedMask_1;
  wire       [7:0]    AlignerPlugin_logic_usedMask_2;
  wire                AlignerPlugin_logic_extractors_0_first;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_usableMask;
  wire       [7:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_2;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_3;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_4;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_5;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_6;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_7;
  reg        [7:0]    _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_slicesOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_3;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_4;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_5;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_6;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_7;
  reg                 AlignerPlugin_logic_extractors_0_redo;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_localMask;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_usageMask;
  reg                 AlignerPlugin_logic_extractors_0_valid;
  reg        [31:0]   AlignerPlugin_logic_extractors_0_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  wire                AlignerPlugin_logic_extractors_0_ctx_trap;
  wire                when_AlignerPlugin_l160;
  wire                AlignerPlugin_logic_extractors_1_first;
  wire       [6:0]    AlignerPlugin_logic_extractors_1_usableMask;
  wire       [6:0]    _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_1;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_2;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_3;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_4;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_5;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_6;
  reg        [6:0]    _zz_AlignerPlugin_logic_extractors_1_slicesOh;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5;
  wire       [6:0]    AlignerPlugin_logic_extractors_1_slicesOh;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_2;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_3;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_4;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_5;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_6;
  reg                 AlignerPlugin_logic_extractors_1_redo;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_localMask;
  wire       [7:0]    AlignerPlugin_logic_extractors_1_usageMask;
  reg                 AlignerPlugin_logic_extractors_1_valid;
  reg        [31:0]   AlignerPlugin_logic_extractors_1_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [3:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [3:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE;
  wire                AlignerPlugin_logic_extractors_1_ctx_trap;
  wire                when_AlignerPlugin_l160_1;
  reg        [9:0]    AlignerPlugin_logic_feeder_harts_0_dopId;
  wire                when_AlignerPlugin_l171;
  wire                AlignerPlugin_logic_feeder_lanes_0_valid;
  wire                AlignerPlugin_logic_feeder_lanes_0_isRvc;
  reg        [31:0]   AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  reg                 AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
  reg        [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
  reg        [14:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
  reg        [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17;
  wire       [12:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21;
  wire       [4:0]    switch_Rvc_l55;
  wire                when_Rvc_l59;
  wire                when_Rvc_l80;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
  wire                when_Rvc_l101;
  wire                when_Rvc_l114;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2;
  reg        [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [1:0]    AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice;
  wire                AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction;
  wire                AlignerPlugin_logic_feeder_lanes_1_valid;
  wire                AlignerPlugin_logic_feeder_lanes_1_isRvc;
  reg        [31:0]   AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
  reg                 AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
  reg        [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
  reg        [14:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
  reg        [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17;
  wire       [12:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21;
  wire       [4:0]    switch_Rvc_l55_1;
  wire                when_Rvc_l59_1;
  wire                when_Rvc_l80_1;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
  wire                when_Rvc_l101_1;
  wire                when_Rvc_l114_1;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2;
  reg        [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3;
  wire       [1:0]    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4;
  wire                _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  wire       [1:0]    AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice;
  wire                AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction;
  reg        [63:0]   AlignerPlugin_logic_buffer_data;
  reg        [3:0]    AlignerPlugin_logic_buffer_mask;
  reg        [3:0]    AlignerPlugin_logic_buffer_last;
  reg        [31:0]   AlignerPlugin_logic_buffer_pc;
  reg                 AlignerPlugin_logic_buffer_trap;
  reg        [9:0]    AlignerPlugin_logic_buffer_hm_Fetch_ID;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3;
  reg        [11:0]   AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY;
  reg        [3:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH;
  reg        [3:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN;
  reg        [31:0]   AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC;
  reg                 AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE;
  wire       [127:0]  _zz_AlignerPlugin_logic_slices_data_0;
  wire                when_AlignerPlugin_l240;
  wire                when_AlignerPlugin_l241;
  wire                when_AlignerPlugin_l241_1;
  wire                AlignerPlugin_logic_buffer_downFire;
  wire       [7:0]    AlignerPlugin_logic_buffer_usedMask;
  wire                AlignerPlugin_logic_buffer_haltUp;
  wire                when_AlignerPlugin_l256;
  wire       [2:0]    _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  wire       [2:0]    _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1;
  wire                when_FpuCsrPlugin_l61;
  wire                LsuPlugin_logic_bus_cmd_valid;
  reg                 LsuPlugin_logic_bus_cmd_ready;
  wire                LsuPlugin_logic_bus_cmd_payload_write;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_address;
  wire       [63:0]   LsuPlugin_logic_bus_cmd_payload_data;
  wire       [1:0]    LsuPlugin_logic_bus_cmd_payload_size;
  wire       [7:0]    LsuPlugin_logic_bus_cmd_payload_mask;
  wire                LsuPlugin_logic_bus_cmd_payload_io;
  wire                LsuPlugin_logic_bus_cmd_payload_fromHart;
  wire       [15:0]   LsuPlugin_logic_bus_cmd_payload_uopId;
  wire                LsuPlugin_logic_bus_rsp_valid;
  wire                LsuPlugin_logic_bus_rsp_payload_error;
  wire       [63:0]   LsuPlugin_logic_bus_rsp_payload_data;
  reg                 LsuPlugin_logic_storeBuffer_push_valid;
  wire       [7:0]    LsuPlugin_logic_storeBuffer_push_payload_slotOh;
  wire       [5:0]    LsuPlugin_logic_storeBuffer_push_payload_tag;
  wire       [31:0]   LsuPlugin_logic_storeBuffer_push_payload_op_address;
  wire       [63:0]   LsuPlugin_logic_storeBuffer_push_payload_op_data;
  wire       [1:0]    LsuPlugin_logic_storeBuffer_push_payload_op_size;
  wire       [11:0]   LsuPlugin_logic_storeBuffer_push_payload_op_storeId;
  wire                LsuPlugin_logic_storeBuffer_pop_valid;
  wire                LsuPlugin_logic_storeBuffer_pop_ready;
  wire       [5:0]    LsuPlugin_logic_storeBuffer_pop_payload_ptr;
  wire       [31:0]   LsuPlugin_logic_storeBuffer_pop_payload_op_address;
  wire       [63:0]   LsuPlugin_logic_storeBuffer_pop_payload_op_data;
  wire       [1:0]    LsuPlugin_logic_storeBuffer_pop_payload_op_size;
  wire       [11:0]   LsuPlugin_logic_storeBuffer_pop_payload_op_storeId;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_ops_pushPtr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_ops_popPtr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_ops_freePtr;
  wire                LsuPlugin_logic_storeBuffer_ops_full;
  wire       [5:0]    LsuPlugin_logic_storeBuffer_ops_occupancy;
  wire       [5:0]    _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address;
  wire       [109:0]  _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1;
  reg                 LsuPlugin_logic_storeBuffer_slots_0_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_0_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_0_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_1_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_1_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_1_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_2_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_2_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_2_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_3_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_3_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_3_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_4_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_4_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_4_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_5_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_5_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_5_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_6_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_6_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_6_tag;
  reg                 LsuPlugin_logic_storeBuffer_slots_7_valid;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_7_ptr;
  reg        [5:0]    LsuPlugin_logic_storeBuffer_slots_7_tag;
  wire                LsuPlugin_logic_storeBuffer_slotsFree;
  wire       [7:0]    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_3;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_4;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_6;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_7;
  reg        [7:0]    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8;
  wire                _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9;
  wire       [7:0]    LsuPlugin_logic_storeBuffer_slotsFreeFirst;
  reg                 LsuPlugin_logic_storeBuffer_holdHart_waitIt;
  wire                when_LsuPlugin_l331;
  reg        [1:0]    LsuPlugin_logic_storeBuffer_waitL1_refill;
  reg                 LsuPlugin_logic_storeBuffer_waitL1_valid;
  wire                when_LsuPlugin_l259;
  wire                LsuPlugin_logic_storeBuffer_empty;
  wire                LsuPlugin_logic_flusher_wantExit;
  reg                 LsuPlugin_logic_flusher_wantStart;
  wire                LsuPlugin_logic_flusher_wantKill;
  reg        [6:0]    LsuPlugin_logic_flusher_cmdCounter;
  wire                LsuPlugin_logic_flusher_inflight;
  reg        [1:0]    LsuPlugin_logic_flusher_waiter;
  wire       [4:0]    LsuPlugin_logic_onAddress0_ls_prefetchOp;
  wire                LsuPlugin_logic_onAddress0_ls_port_valid;
  wire                LsuPlugin_logic_onAddress0_ls_port_ready;
  reg        [2:0]    LsuPlugin_logic_onAddress0_ls_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_ls_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_ls_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_ls_port_payload_storeId;
  reg        [11:0]   LsuPlugin_logic_onAddress0_ls_storeId;
  wire                LsuPlugin_logic_onAddress0_ls_port_fire;
  wire                LsuPlugin_logic_onAddress0_flush_port_valid;
  wire                LsuPlugin_logic_onAddress0_flush_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_flush_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_flush_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_flush_port_payload_storeId;
  wire                LsuPlugin_logic_onAddress0_flush_port_fire;
  wire                LsuPlugin_logic_onAddress0_sb_isHead;
  wire                LsuPlugin_logic_onAddress0_sb_flush;
  wire                LsuPlugin_logic_onAddress0_sb_port_valid;
  wire                LsuPlugin_logic_onAddress0_sb_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_sb_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_sb_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_sb_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_sb_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_sb_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_sb_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_sb_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_sb_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_sb_port_payload_storeId;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_valid;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_fromHp_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_fromHp_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_fromHp_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_fromHp_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_fromHp_port_payload_storeId;
  reg        [7:0]    _zz_execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                when_LsuPlugin_l546;
  wire                when_LsuPlugin_l546_1;
  wire       [31:0]   LsuPlugin_logic_onPma_cached_cmd_address;
  wire       [0:0]    LsuPlugin_logic_onPma_cached_cmd_op;
  wire                LsuPlugin_logic_onPma_cached_rsp_fault;
  wire                LsuPlugin_logic_onPma_cached_rsp_io;
  wire       [31:0]   LsuPlugin_logic_onPma_io_cmd_address;
  wire       [1:0]    LsuPlugin_logic_onPma_io_cmd_size;
  wire       [0:0]    LsuPlugin_logic_onPma_io_cmd_op;
  wire                LsuPlugin_logic_onPma_io_rsp_fault;
  wire                LsuPlugin_logic_onPma_io_rsp_io;
  wire                when_LsuPlugin_l569;
  wire                LsuPlugin_logic_onPma_addressExtension;
  reg                 LsuPlugin_logic_onCtrl_lsuTrap;
  reg        [63:0]   LsuPlugin_logic_onCtrl_writeData;
  wire                LsuPlugin_logic_onCtrl_scMiss;
  reg                 LsuPlugin_logic_onCtrl_io_tooEarly;
  reg                 LsuPlugin_logic_onCtrl_io_allowIt;
  wire                when_LsuPlugin_l597;
  wire                LsuPlugin_logic_onCtrl_io_doIt;
  reg                 LsuPlugin_logic_onCtrl_io_doItReg;
  reg                 LsuPlugin_logic_onCtrl_io_cmdSent;
  wire                LsuPlugin_logic_bus_cmd_fire;
  wire                when_LsuPlugin_l601;
  wire                LsuPlugin_logic_bus_rsp_toStream_valid;
  wire                LsuPlugin_logic_bus_rsp_toStream_ready;
  wire                LsuPlugin_logic_bus_rsp_toStream_payload_error;
  wire       [63:0]   LsuPlugin_logic_bus_rsp_toStream_payload_data;
  wire                LsuPlugin_logic_onCtrl_io_rsp_valid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_ready;
  wire                LsuPlugin_logic_onCtrl_io_rsp_payload_error;
  wire       [63:0]   LsuPlugin_logic_onCtrl_io_rsp_payload_data;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rValid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_fire;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rData_error;
  reg        [63:0]   LsuPlugin_logic_bus_rsp_toStream_rData_data;
  wire                LsuPlugin_logic_onCtrl_io_freezeIt;
  wire       [63:0]   LsuPlugin_logic_onCtrl_loadData_input;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_0;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_1;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_2;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_3;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_4;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_5;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_6;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_7;
  reg        [63:0]   LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
  wire       [63:0]   LsuPlugin_logic_onCtrl_storeData_mapping_3_1;
  reg        [63:0]   _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_srcBuffer;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire                LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                LsuPlugin_logic_onCtrl_rva_alu_unsigned;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire                LsuPlugin_logic_onCtrl_rva_alu_less;
  wire                LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire       [2:0]    switch_Misc_l245;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_alu_raw;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_result;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_aluBuffer;
  wire                LsuPlugin_logic_onCtrl_rva_delay_0;
  wire                LsuPlugin_logic_onCtrl_rva_delay_1;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  wire                LsuPlugin_logic_onCtrl_rva_freezeIt;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_capture;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_lrsc_address;
  wire                when_LsuPlugin_l686;
  reg        [5:0]    LsuPlugin_logic_onCtrl_rva_lrsc_age;
  wire                when_LsuPlugin_l698;
  wire                when_LsuPlugin_l705;
  wire                when_LsuPlugin_l709;
  wire       [5:0]    LsuPlugin_logic_onCtrl_wb_tag;
  wire       [7:0]    LsuPlugin_logic_onCtrl_wb_hits;
  wire                LsuPlugin_logic_onCtrl_wb_hit;
  wire                LsuPlugin_logic_onCtrl_wb_compatibleOp;
  wire                LsuPlugin_logic_onCtrl_wb_notFull;
  wire                LsuPlugin_logic_onCtrl_wb_allowed;
  wire       [7:0]    LsuPlugin_logic_onCtrl_wb_slotOh;
  wire                LsuPlugin_logic_onCtrl_wb_loadHazard;
  wire                LsuPlugin_logic_onCtrl_wb_selfHazard;
  wire                LsuPlugin_logic_onCtrl_traps_accessFault;
  wire                LsuPlugin_logic_onCtrl_traps_l1Failed;
  wire                when_LsuPlugin_l759;
  wire                LsuPlugin_logic_onCtrl_traps_pmaFault;
  wire                when_LsuPlugin_l810;
  wire                when_LsuPlugin_l837;
  wire                LsuPlugin_logic_onCtrl_fenceTrap_valid;
  wire                when_LsuPlugin_l865;
  wire                when_LsuPlugin_l873;
  wire                when_LsuPlugin_l876;
  wire                LsuPlugin_logic_onCtrl_mmuNeeded;
  wire                when_LsuPlugin_l905;
  wire                when_LsuPlugin_l910;
  wire                when_LsuPlugin_l913;
  wire                when_LsuPlugin_l263;
  wire                when_LsuPlugin_l918;
  wire                when_LsuPlugin_l918_1;
  wire                when_LsuPlugin_l918_2;
  wire                when_LsuPlugin_l918_3;
  wire                when_LsuPlugin_l918_4;
  wire                when_LsuPlugin_l918_5;
  wire                when_LsuPlugin_l918_6;
  wire                when_LsuPlugin_l918_7;
  reg        [1:0]    LsuPlugin_logic_onCtrl_hartRegulation_refill;
  reg                 LsuPlugin_logic_onCtrl_hartRegulation_valid;
  wire                when_LsuPlugin_l259_1;
  wire                when_LsuPlugin_l949;
  wire                when_LsuPlugin_l263_1;
  wire                LsuPlugin_logic_onCtrl_commitProbeReq;
  reg                 LsuPlugin_logic_onCtrl_commitProbeToken;
  wire                when_LsuPlugin_l974;
  wire                when_LsuPlugin_l982;
  wire                LsuPlugin_logic_onWb_storeFire;
  wire                LsuPlugin_logic_onWb_storeBroadcast;
  wire                when_StageLink_l71_1;
  wire                when_StageLink_l71_2;
  wire                FpuPackerPlugin_logic_flagsWb_flags_NX;
  wire                FpuPackerPlugin_logic_flagsWb_flags_UF;
  wire                FpuPackerPlugin_logic_flagsWb_flags_OF;
  wire                FpuPackerPlugin_logic_flagsWb_flags_DZ;
  wire                FpuPackerPlugin_logic_flagsWb_flags_NV;
  wire       [4:0]    FpuPackerPlugin_logic_flagsWb_ats;
  wire                FpuPackerPlugin_wb_at_2_valid;
  wire       [63:0]   FpuPackerPlugin_wb_at_2_payload;
  wire                FpuPackerPlugin_wb_at_5_valid;
  wire       [63:0]   FpuPackerPlugin_wb_at_5_payload;
  wire                FpuPackerPlugin_wb_at_3_valid;
  wire       [63:0]   FpuPackerPlugin_wb_at_3_payload;
  wire                FpuPackerPlugin_wb_at_6_valid;
  wire       [63:0]   FpuPackerPlugin_wb_at_6_payload;
  wire                FpuPackerPlugin_wb_at_9_valid;
  wire       [63:0]   FpuPackerPlugin_wb_at_9_payload;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_0_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_0_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_0_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_0_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_0_mantissa;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_1_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_1_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_1_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_1_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_1_mantissa;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_2_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_2_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_2_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_2_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_2_mantissa;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_3_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_3_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_3_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_3_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_3_mantissa;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_4_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_4_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_4_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_4_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_4_mantissa;
  wire       [1:0]    FpuPackerPlugin_logic_s0_remapped_5_mode;
  wire                FpuPackerPlugin_logic_s0_remapped_5_quiet;
  wire                FpuPackerPlugin_logic_s0_remapped_5_sign;
  wire       [12:0]   FpuPackerPlugin_logic_s0_remapped_5_exponent;
  wire       [53:0]   FpuPackerPlugin_logic_s0_remapped_5_mantissa;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid_1;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid_2;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid_3;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid_4;
  wire                _zz_FpuPackerPlugin_logic_pip_node_0_valid_5;
  wire       [5:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet;
  wire       [1:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode;
  wire       [70:0]   _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1;
  wire       [1:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1;
  wire       [0:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT;
  wire       [0:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1;
  wire       [2:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE;
  wire       [2:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1;
  wire       [4:0]    _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX;
  wire       [2:0]    _zz_49;
  wire       [2:0]    _zz_50;
  wire       [2:0]    _zz_51;
  wire       [2:0]    _zz_52;
  wire       [2:0]    _zz_53;
  wire       [2:0]    _zz_54;
  wire       [2:0]    _zz_55;
  wire       [2:0]    _zz_56;
  wire       [12:0]   _zz_when_AFix_l1168_1;
  reg        [12:0]   _zz_FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE;
  wire                when_AFix_l1168_1;
  reg        [5:0]    _zz_FpuPackerPlugin_logic_s1_subnormal_manShift;
  wire                when_UInt_l119_1;
  reg        [5:0]    FpuPackerPlugin_logic_s1_subnormal_manShift;
  wire       [54:0]   _zz_when_Utils_l1585_15;
  reg                 _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1;
  wire                when_Utils_l1585_7;
  wire                when_Utils_l1585_8;
  wire                when_Utils_l1585_9;
  wire                when_Utils_l1585_10;
  wire                when_Utils_l1585_11;
  wire                when_Utils_l1585_12;
  reg        [53:0]   FpuPackerPlugin_logic_s1_subnormal_manShifter;
  reg        [1:0]    FpuPackerPlugin_logic_s1_subnormal_counter;
  wire                FpuPackerPlugin_logic_s1_subnormal_freezeIt;
  wire                when_FpuPackerPlugin_l134;
  reg                 _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR;
  wire       [29:0]   FpuPackerPlugin_logic_s1_incrBy;
  wire       [52:0]   FpuPackerPlugin_logic_s1_manIncrWithCarry;
  wire                FpuPackerPlugin_logic_s1_MAN_CARRY;
  wire       [51:0]   FpuPackerPlugin_logic_s1_MAN_INCR;
  wire       [1:0]    FpuPackerPlugin_logic_s2_tinyRound;
  reg                 _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr;
  wire                FpuPackerPlugin_logic_s2_tinyRoundingIncr;
  wire                FpuPackerPlugin_logic_s2_tinyOverflow;
  reg                 FpuPackerPlugin_logic_s2_expSet;
  reg                 FpuPackerPlugin_logic_s2_expZero;
  reg                 FpuPackerPlugin_logic_s2_expMax;
  reg                 FpuPackerPlugin_logic_s2_manZero;
  reg                 FpuPackerPlugin_logic_s2_manSet;
  reg                 FpuPackerPlugin_logic_s2_manOne;
  reg                 FpuPackerPlugin_logic_s2_manQuiet;
  reg                 FpuPackerPlugin_logic_s2_positive;
  reg                 FpuPackerPlugin_logic_s2_nx;
  reg                 FpuPackerPlugin_logic_s2_of;
  reg                 FpuPackerPlugin_logic_s2_uf;
  wire                when_FpuPackerPlugin_l208;
  wire                when_FpuPackerPlugin_l210;
  reg                 when_FpuPackerPlugin_l224;
  reg                 _zz_when_FpuPackerPlugin_l241;
  wire                when_FpuPackerPlugin_l241;
  wire                FpuPackerPlugin_logic_s2_fwb_flags_NX;
  wire                FpuPackerPlugin_logic_s2_fwb_flags_UF;
  wire                FpuPackerPlugin_logic_s2_fwb_flags_OF;
  wire                FpuPackerPlugin_logic_s2_fwb_flags_DZ;
  wire                FpuPackerPlugin_logic_s2_fwb_flags_NV;
  reg        [63:0]   FpuPackerPlugin_logic_s2_fwb_value;
  wire                FpuPackerPlugin_logic_s2_fpWriter_valid;
  wire       [15:0]   FpuPackerPlugin_logic_s2_fpWriter_payload_uopId;
  wire       [63:0]   FpuPackerPlugin_logic_s2_fpWriter_payload_data;
  wire                when_Misc_l22;
  wire                when_Misc_l22_1;
  wire                when_Misc_l22_2;
  wire                when_Misc_l22_3;
  wire                when_Misc_l22_4;
  wire                when_Misc_l22_5;
  wire                when_Misc_l22_6;
  wire                when_Misc_l22_7;
  wire                when_Misc_l22_8;
  wire                when_FpuPackerPlugin_l309;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [1:0]    CsrRamPlugin_setup_initPort_address;
  wire       [31:0]   CsrRamPlugin_setup_initPort_data;
  wire                early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l245_1;
  reg                 _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                early0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early0_BranchPlugin_logic_jumpLogic_needFix;
  wire                early0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_history_slice;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l213;
  wire                when_BranchPlugin_l213_1;
  wire                when_BranchPlugin_l213_2;
  wire                when_BranchPlugin_l218;
  wire                early0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                early1_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l245_2;
  reg                 _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
  reg                 _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  wire                early1_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early1_BranchPlugin_logic_jumpLogic_needFix;
  wire                early1_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    early1_BranchPlugin_logic_jumpLogic_history_slice;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l213_3;
  wire                when_BranchPlugin_l213_4;
  wire                when_BranchPlugin_l213_5;
  wire                when_BranchPlugin_l218_1;
  wire                early1_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early1_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early1_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                PmpPlugin_logic_isMachine;
  wire                PmpPlugin_logic_instructionShouldHit;
  wire                PmpPlugin_logic_dataShouldHit;
  wire                FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   FetchL1Plugin_logic_pmpPort_logic_torCmpAddress;
  wire                LsuPlugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   LsuPlugin_logic_pmpPort_logic_torCmpAddress;
  wire                LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid;
  wire                LsuCachelessWishbonePlugin_logic_bridge_cmdStage_ready;
  wire                LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_write;
  wire       [31:0]   LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_address;
  wire       [63:0]   LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_data;
  wire       [1:0]    LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_size;
  wire       [7:0]    LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_mask;
  wire                LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_io;
  wire                LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_fromHart;
  wire       [15:0]   LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_uopId;
  reg                 LsuPlugin_logic_bus_cmd_rValid;
  reg                 LsuPlugin_logic_bus_cmd_rData_write;
  reg        [31:0]   LsuPlugin_logic_bus_cmd_rData_address;
  reg        [63:0]   LsuPlugin_logic_bus_cmd_rData_data;
  reg        [1:0]    LsuPlugin_logic_bus_cmd_rData_size;
  reg        [7:0]    LsuPlugin_logic_bus_cmd_rData_mask;
  reg                 LsuPlugin_logic_bus_cmd_rData_io;
  reg                 LsuPlugin_logic_bus_cmd_rData_fromHart;
  reg        [15:0]   LsuPlugin_logic_bus_cmd_rData_uopId;
  wire                when_Stream_l477_2;
  wire                LsuPlugin_logic_commitProbe_takeWhen_valid;
  wire       [31:0]   LsuPlugin_logic_commitProbe_takeWhen_payload_pc;
  wire       [31:0]   LsuPlugin_logic_commitProbe_takeWhen_payload_address;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_load;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_store;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_trap;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_io;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_prefetchFailed;
  wire                LsuPlugin_logic_commitProbe_takeWhen_payload_miss;
  wire                when_Prefetcher_l155;
  wire       [3:0]    _zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT;
  wire                PrefetcherRptPlugin_logic_onCtrl_unfiltred_valid;
  wire                PrefetcherRptPlugin_logic_onCtrl_unfiltred_ready;
  wire       [31:0]   PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_address;
  wire                PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_unique;
  wire       [2:0]    PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_from;
  wire       [2:0]    PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to;
  wire       [11:0]   PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride;
  reg        [4:0]    PrefetcherRptPlugin_logic_onCtrl_add;
  reg        [4:0]    PrefetcherRptPlugin_logic_onCtrl_sub;
  wire       [5:0]    _zz_when_UInt_l128;
  reg        [4:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_score;
  wire                when_UInt_l128;
  wire       [5:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_score_1;
  reg        [4:0]    PrefetcherRptPlugin_logic_onCtrl_score;
  wire                when_UInt_l119_2;
  wire       [3:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed;
  reg        [2:0]    PrefetcherRptPlugin_logic_onCtrl_advanceSubed;
  wire                when_UInt_l128_1;
  wire       [5:0]    _zz_when_UInt_l128_1;
  reg        [4:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_advanceAllowed;
  wire                when_UInt_l128_2;
  wire       [4:0]    PrefetcherRptPlugin_logic_onCtrl_advanceAllowed;
  reg                 PrefetcherRptPlugin_logic_onCtrl_orderAsk;
  wire                PrefetcherRptPlugin_logic_onCtrl_unfiltred_fire;
  wire       [2:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to;
  wire       [6:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride;
  wire       [7:0]    _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1;
  wire                when_Prefetcher_l196;
  wire                when_Prefetcher_l197;
  wire                when_Prefetcher_l198;
  wire                when_Prefetcher_l208;
  wire                when_Prefetcher_l216;
  wire       [31:0]   LsuPlugin_pmaBuilder_l1_addressBits;
  wire       [0:0]    LsuPlugin_pmaBuilder_l1_argsBits;
  wire                _zz_LsuPlugin_logic_onPma_cached_rsp_io;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_io_addressBits;
  wire       [2:0]    LsuPlugin_pmaBuilder_io_argsBits;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_hit;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_fault;
  wire                _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  wire                _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX;
  wire                _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1;
  wire                _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_0_UF;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_0_OF;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_0_DZ;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NV;
  wire                execute_lane0_ctrls_7_upIsCancel;
  wire                execute_lane0_ctrls_7_downIsCancel;
  wire                execute_lane0_ctrls_5_upIsCancel;
  wire                execute_lane0_ctrls_5_downIsCancel;
  wire                execute_lane0_ctrls_8_upIsCancel;
  wire                execute_lane0_ctrls_8_downIsCancel;
  wire                execute_lane0_ctrls_11_upIsCancel;
  wire                execute_lane0_ctrls_11_downIsCancel;
  wire                _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_1_UF;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_1_OF;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_1_DZ;
  wire                FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NV;
  wire                FpuFlagsWritebackPlugin_logic_flagsOr_NX;
  wire                FpuFlagsWritebackPlugin_logic_flagsOr_UF;
  wire                FpuFlagsWritebackPlugin_logic_flagsOr_OF;
  wire                FpuFlagsWritebackPlugin_logic_flagsOr_DZ;
  wire                FpuFlagsWritebackPlugin_logic_flagsOr_NV;
  wire                CsrRamPlugin_csrMapper_read_valid;
  wire                CsrRamPlugin_csrMapper_read_ready;
  wire       [1:0]    CsrRamPlugin_csrMapper_read_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_read_data;
  wire                CsrRamPlugin_csrMapper_write_valid;
  wire                CsrRamPlugin_csrMapper_write_ready;
  wire       [1:0]    CsrRamPlugin_csrMapper_write_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_write_data;
  wire                late0_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l245_3;
  reg                 _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                late0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                late0_BranchPlugin_logic_jumpLogic_needFix;
  wire                late0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_history_slice;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l213_6;
  wire                when_BranchPlugin_l213_7;
  wire                when_BranchPlugin_l213_8;
  wire                when_BranchPlugin_l218_2;
  wire                late0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                late0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                late0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_valid;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                late1_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l245_4;
  reg                 _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  reg                 _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  wire                late1_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                late1_BranchPlugin_logic_jumpLogic_needFix;
  wire                late1_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_history_slice;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l213_9;
  wire                when_BranchPlugin_l213_10;
  wire                when_BranchPlugin_l213_11;
  wire                when_BranchPlugin_l218_3;
  wire                late1_BranchPlugin_logic_jumpLogic_rdLink;
  wire                late1_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                late1_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_valid;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                execute_lane0_ctrls_10_upIsCancel;
  wire                execute_lane0_ctrls_10_downIsCancel;
  wire       [1:0]    CsrRamPlugin_csrMapper_ramAddress;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress;
  reg                 CsrRamPlugin_csrMapper_withRead;
  wire                when_CsrRamPlugin_l85;
  reg                 CsrRamPlugin_csrMapper_doWrite;
  reg                 CsrRamPlugin_csrMapper_fired;
  wire                when_CsrRamPlugin_l92;
  wire                when_CsrRamPlugin_l96;
  wire                LearnPlugin_logic_learn_valid;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcTarget;
  wire                LearnPlugin_logic_learn_payload_taken;
  wire                LearnPlugin_logic_learn_payload_isBranch;
  wire                LearnPlugin_logic_learn_payload_isPush;
  wire                LearnPlugin_logic_learn_payload_isPop;
  wire                LearnPlugin_logic_learn_payload_wasWrong;
  wire                LearnPlugin_logic_learn_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_learn_payload_history;
  wire       [15:0]   LearnPlugin_logic_learn_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                LearnPlugin_logic_buffered_0_valid;
  wire                LearnPlugin_logic_buffered_0_ready;
  wire       [31:0]   LearnPlugin_logic_buffered_0_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_buffered_0_payload_pcTarget;
  wire                LearnPlugin_logic_buffered_0_payload_taken;
  wire                LearnPlugin_logic_buffered_0_payload_isBranch;
  wire                LearnPlugin_logic_buffered_0_payload_isPush;
  wire                LearnPlugin_logic_buffered_0_payload_isPop;
  wire                LearnPlugin_logic_buffered_0_payload_wasWrong;
  wire                LearnPlugin_logic_buffered_0_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_buffered_0_payload_history;
  wire       [15:0]   LearnPlugin_logic_buffered_0_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rValid;
  reg        [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  reg        [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_history;
  reg        [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                when_Stream_l477_3;
  wire                LearnPlugin_logic_buffered_1_valid;
  wire                LearnPlugin_logic_buffered_1_ready;
  wire       [31:0]   LearnPlugin_logic_buffered_1_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_buffered_1_payload_pcTarget;
  wire                LearnPlugin_logic_buffered_1_payload_taken;
  wire                LearnPlugin_logic_buffered_1_payload_isBranch;
  wire                LearnPlugin_logic_buffered_1_payload_isPush;
  wire                LearnPlugin_logic_buffered_1_payload_isPop;
  wire                LearnPlugin_logic_buffered_1_payload_wasWrong;
  wire                LearnPlugin_logic_buffered_1_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_buffered_1_payload_history;
  wire       [15:0]   LearnPlugin_logic_buffered_1_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rValid;
  reg        [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  reg        [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_history;
  reg        [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                when_Stream_l477_4;
  wire                LearnPlugin_logic_arbitrated_valid;
  wire                LearnPlugin_logic_arbitrated_ready;
  wire       [31:0]   LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_arbitrated_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_payload_taken;
  wire                LearnPlugin_logic_arbitrated_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                LearnPlugin_logic_arbitrated_toFlow_valid;
  wire       [31:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_toFlow_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  reg        [15:0]   DecoderPlugin_logic_harts_0_uopId;
  wire                when_DecoderPlugin_l143;
  wire       [0:0]    DecoderPlugin_logic_interrupt_async;
  wire                when_DecoderPlugin_l151;
  reg        [0:0]    DecoderPlugin_logic_interrupt_buffered;
  wire                _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire                _zz_decode_ctrls_1_down_RD_RFID_0;
  wire                _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_0_fp_instRm;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_0_fp_rm;
  wire                DecoderPlugin_logic_laneLogic_0_fp_triggered;
  wire                DecoderPlugin_logic_laneLogic_0_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  wire       [31:0]   DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50_2;
  wire                when_DecoderPlugin_l229;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  wire                when_DecoderPlugin_l247;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_uopIdBase;
  wire                _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1;
  wire                _zz_decode_ctrls_1_down_RD_RFID_1;
  wire                _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_1_fp_instRm;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_1_fp_rm;
  wire                DecoderPlugin_logic_laneLogic_1_fp_triggered;
  wire                DecoderPlugin_logic_laneLogic_1_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_1_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception;
  wire       [31:0]   DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_code;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1;
  wire                DecoderPlugin_logic_laneLogic_1_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_1_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit;
  reg                 decode_ctrls_1_up_LANE_SEL_1_regNext;
  wire                when_CtrlLaneApi_l50_3;
  wire                when_DecoderPlugin_l229_1;
  wire                DecoderPlugin_logic_laneLogic_1_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_1_flushPort_payload_self;
  wire                when_DecoderPlugin_l247_1;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_uopIdBase;
  reg                 DispatchPlugin_logic_slots_0_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_laneLayerHits;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_uop;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  reg        [11:0]   DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_hm_PC;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_TRAP;
  reg        [15:0]   DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS1_RFID;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS2_RFID;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_RD_RFID;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RS3_ENABLE;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS3_RFID;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS3_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_valid;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_uop;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_fire;
  wire                DispatchPlugin_logic_candidates_0_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_0_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_0_reservationHazards;
  wire                DispatchPlugin_logic_candidates_0_flushHazards;
  wire                DispatchPlugin_logic_candidates_0_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_age;
  wire                DispatchPlugin_logic_candidates_0_moving;
  wire                DispatchPlugin_logic_candidates_1_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_uop;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_fire;
  wire                DispatchPlugin_logic_candidates_1_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_reservationHazards;
  wire                DispatchPlugin_logic_candidates_1_flushHazards;
  wire                DispatchPlugin_logic_candidates_1_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_age;
  wire                DispatchPlugin_logic_candidates_1_moving;
  wire                DispatchPlugin_logic_candidates_2_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_uop;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_fire;
  wire                DispatchPlugin_logic_candidates_2_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_reservationHazards;
  wire                DispatchPlugin_logic_candidates_2_flushHazards;
  wire                DispatchPlugin_logic_candidates_2_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_age;
  wire                DispatchPlugin_logic_candidates_2_moving;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_2_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_2_hazard;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_0_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_2_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_0_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_2_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_0_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_2_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_3_hit;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_oldersHazard;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_1_oldersHazard;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_2_oldersHazard;
  wire       [0:0]    DispatchPlugin_logic_fenceChecker_olderInflights;
  wire                DispatchPlugin_logic_feeds_0_sending;
  reg                 DispatchPlugin_logic_feeds_0_sent;
  wire                when_DispatchPlugin_l368;
  wire                DispatchPlugin_logic_feeds_1_sending;
  reg                 DispatchPlugin_logic_feeds_1_sent;
  wire                when_DispatchPlugin_l368_1;
  wire                when_DispatchPlugin_l378;
  wire       [1:0]    _zz_GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_1;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_2;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_3;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l119;
  wire                when_GSharePlugin_l119_1;
  wire                when_GSharePlugin_l119_2;
  wire                when_GSharePlugin_l119_3;
  wire       [11:0]   BtbPlugin_logic_onLearn_hash;
  wire       [22:0]   FpuUnpack_RS1_f32_mantissa;
  wire       [7:0]    FpuUnpack_RS1_f32_exponent;
  wire                FpuUnpack_RS1_f32_sign;
  wire       [51:0]   FpuUnpack_RS1_f64_mantissa;
  wire       [10:0]   FpuUnpack_RS1_f64_exponent;
  wire                FpuUnpack_RS1_f64_sign;
  reg                 FpuUnpack_RS1_manZero;
  reg                 FpuUnpack_RS1_expZero;
  reg                 FpuUnpack_RS1_expOne;
  reg        [11:0]   FpuUnpack_RS1_recodedExpSub;
  wire                when_Misc_l22_9;
  wire       [1:0]    switch_Misc_l245_5;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1;
  reg        [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2;
  wire                FpuUnpack_RS1_normalizer_unpackerSel;
  wire                FpuUnpack_RS1_normalizer_valid;
  reg                 FpuUnpack_RS1_normalizer_validReg;
  wire                when_FpuUnpackerPlugin_l234;
  reg                 FpuUnpack_RS1_normalizer_asked;
  wire                when_FpuUnpackerPlugin_l235;
  reg                 FpuUnpack_RS1_normalizer_served;
  wire                when_FpuUnpackerPlugin_l236;
  reg        [11:0]   FpuUnpack_RS1_normalizer_exponent;
  reg        [51:0]   FpuUnpack_RS1_normalizer_mantissa;
  wire                when_FpuUnpackerPlugin_l243;
  wire                when_FpuUnpackerPlugin_l251;
  wire                FpuUnpack_RS1_normalizer_freezeIt;
  wire       [22:0]   FpuUnpack_RS2_f32_mantissa;
  wire       [7:0]    FpuUnpack_RS2_f32_exponent;
  wire                FpuUnpack_RS2_f32_sign;
  wire       [51:0]   FpuUnpack_RS2_f64_mantissa;
  wire       [10:0]   FpuUnpack_RS2_f64_exponent;
  wire                FpuUnpack_RS2_f64_sign;
  reg                 FpuUnpack_RS2_manZero;
  reg                 FpuUnpack_RS2_expZero;
  reg                 FpuUnpack_RS2_expOne;
  reg        [11:0]   FpuUnpack_RS2_recodedExpSub;
  wire                when_Misc_l22_10;
  wire       [1:0]    switch_Misc_l245_6;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1;
  reg        [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2;
  wire                FpuUnpack_RS2_normalizer_unpackerSel;
  wire                FpuUnpack_RS2_normalizer_valid;
  reg                 FpuUnpack_RS2_normalizer_validReg;
  wire                when_FpuUnpackerPlugin_l234_1;
  reg                 FpuUnpack_RS2_normalizer_asked;
  wire                when_FpuUnpackerPlugin_l235_1;
  reg                 FpuUnpack_RS2_normalizer_served;
  wire                when_FpuUnpackerPlugin_l236_1;
  reg        [11:0]   FpuUnpack_RS2_normalizer_exponent;
  reg        [51:0]   FpuUnpack_RS2_normalizer_mantissa;
  wire                when_FpuUnpackerPlugin_l243_1;
  wire                when_FpuUnpackerPlugin_l251_1;
  wire                FpuUnpack_RS2_normalizer_freezeIt;
  wire       [22:0]   FpuUnpack_RS3_f32_mantissa;
  wire       [7:0]    FpuUnpack_RS3_f32_exponent;
  wire                FpuUnpack_RS3_f32_sign;
  wire       [51:0]   FpuUnpack_RS3_f64_mantissa;
  wire       [10:0]   FpuUnpack_RS3_f64_exponent;
  wire                FpuUnpack_RS3_f64_sign;
  reg                 FpuUnpack_RS3_manZero;
  reg                 FpuUnpack_RS3_expZero;
  reg                 FpuUnpack_RS3_expOne;
  reg        [11:0]   FpuUnpack_RS3_recodedExpSub;
  wire                when_Misc_l22_11;
  wire       [1:0]    switch_Misc_l245_7;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode;
  wire       [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1;
  reg        [1:0]    _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2;
  wire                FpuUnpack_RS3_normalizer_unpackerSel;
  wire                FpuUnpack_RS3_normalizer_valid;
  reg                 FpuUnpack_RS3_normalizer_validReg;
  wire                when_FpuUnpackerPlugin_l234_2;
  reg                 FpuUnpack_RS3_normalizer_asked;
  wire                when_FpuUnpackerPlugin_l235_2;
  reg                 FpuUnpack_RS3_normalizer_served;
  wire                when_FpuUnpackerPlugin_l236_2;
  reg        [11:0]   FpuUnpack_RS3_normalizer_exponent;
  reg        [51:0]   FpuUnpack_RS3_normalizer_mantissa;
  wire                when_FpuUnpackerPlugin_l243_2;
  wire                when_FpuUnpackerPlugin_l251_2;
  wire                FpuUnpack_RS3_normalizer_freezeIt;
  wire                FpuUnpackerPlugin_logic_unpackDone;
  wire                FpuUnpackerPlugin_logic_onCvt_rs1Zero;
  reg                 FpuUnpackerPlugin_logic_onCvt_asked;
  reg                 FpuUnpackerPlugin_logic_onCvt_served;
  reg        [5:0]    FpuUnpackerPlugin_logic_onCvt_fsmResult_shift;
  reg        [51:0]   FpuUnpackerPlugin_logic_onCvt_fsmResult_data;
  wire                FpuUnpackerPlugin_logic_onCvt_freezeIt;
  wire       [4:0]    _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [0:0]    lane0_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire                lane0_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane0_integer_WriteBackPlugin_logic_write_port_address;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  wire       [1:0]    lane1_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane1_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [1:0]    lane1_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane1_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire                lane1_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane1_integer_WriteBackPlugin_logic_write_port_address;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_write_port_uopId;
  wire       [0:0]    lane0_float_WriteBackPlugin_logic_stages_0_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane0_float_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [2:0]    lane0_float_WriteBackPlugin_logic_stages_1_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_1_muxed;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_1_merged;
  wire                lane0_float_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [0:0]    lane0_float_WriteBackPlugin_logic_stages_2_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_2_muxed;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_2_merged;
  wire                lane0_float_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire       [0:0]    lane0_float_WriteBackPlugin_logic_stages_3_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_3_muxed;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_3_merged;
  wire                lane0_float_WriteBackPlugin_logic_stages_3_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_3_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_3_write_payload_data;
  wire       [0:0]    lane0_float_WriteBackPlugin_logic_stages_4_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_4_muxed;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_4_merged;
  wire                lane0_float_WriteBackPlugin_logic_stages_4_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_4_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_4_write_payload_data;
  wire       [0:0]    lane0_float_WriteBackPlugin_logic_stages_5_hits;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_5_muxed;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_5_merged;
  wire                lane0_float_WriteBackPlugin_logic_stages_5_write_valid;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_stages_5_write_payload_uopId;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_stages_5_write_payload_data;
  wire                lane0_float_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane0_float_WriteBackPlugin_logic_write_port_address;
  wire       [63:0]   lane0_float_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane0_float_WriteBackPlugin_logic_write_port_uopId;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_7;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_8;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_9;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_10;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_11;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_12;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_13;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_14;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_15;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1;
  wire                _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_7;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_8;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_9;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_10;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_11;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_12;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_13;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_14;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_15;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1;
  wire                _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1;
  reg        [9:0]    FpuClassPlugin_logic_onWb_fclassResult;
  wire       [10:0]   FpuClassPlugin_logic_onWb_expSubnormal;
  wire                FpuCmpPlugin_logic_onCmp_signalQuiet;
  wire                FpuCmpPlugin_logic_onCmp_rs1NanNv;
  wire                FpuCmpPlugin_logic_onCmp_rs2NanNv;
  reg                 FpuCmpPlugin_logic_onCmp_rs1AbsSmaller;
  wire                when_FpuCmpPlugin_l110;
  wire                when_FpuCmpPlugin_l111;
  wire                when_FpuCmpPlugin_l112;
  wire                when_FpuCmpPlugin_l113;
  wire                when_FpuCmpPlugin_l114;
  wire       [1:0]    switch_Misc_l245_8;
  reg                 FpuCmpPlugin_logic_onCmp_rs1Smaller;
  wire                when_FpuCmpPlugin_l124;
  reg                 FpuCmpPlugin_logic_onFloatWb_doNan;
  wire                when_Misc_l22_12;
  wire                when_Misc_l22_13;
  wire                when_Misc_l22_14;
  wire                when_Misc_l22_15;
  wire                when_FpuCmpPlugin_l149;
  wire                when_FpuCmpPlugin_l153;
  wire                when_Misc_l22_16;
  wire       [11:0]   _zz_when_UInt_l119;
  reg        [5:0]    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  wire                when_UInt_l119_3;
  wire       [53:0]   _zz_when_Utils_l1585_16;
  wire       [3:0]    _zz_when_Utils_l1585_17;
  reg                 _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1;
  wire                when_Utils_l1585_13;
  wire                when_Utils_l1585_14;
  wire                when_Utils_l1585_15;
  wire                when_Utils_l1585_16;
  wire                FpuF2iPlugin_logic_onShift_signed;
  wire       [5:0]    _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6;
  reg                 _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  wire                when_Utils_l1585_17;
  wire                when_Utils_l1585_18;
  wire                when_Utils_l1585_19;
  wire                when_Utils_l1585_20;
  wire                when_Utils_l1585_21;
  wire                when_Utils_l1585_22;
  wire       [31:0]   FpuF2iPlugin_logic_onShift_high;
  wire       [21:0]   FpuF2iPlugin_logic_onShift_low;
  wire       [31:0]   FpuF2iPlugin_logic_onShift_unsigned;
  wire       [1:0]    FpuF2iPlugin_logic_onShift_round;
  reg                 _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0;
  wire                FpuF2iPlugin_logic_onResult_signed;
  wire                FpuF2iPlugin_logic_onResult_i64;
  wire       [31:0]   FpuF2iPlugin_logic_onResult_high;
  wire       [21:0]   FpuF2iPlugin_logic_onResult_low;
  wire       [31:0]   FpuF2iPlugin_logic_onResult_unsigned;
  wire       [1:0]    FpuF2iPlugin_logic_onResult_round;
  reg                 FpuF2iPlugin_logic_onResult_halfRater_firstCycle;
  wire                FpuF2iPlugin_logic_onResult_halfRater_freezeIt;
  reg        [31:0]   FpuF2iPlugin_logic_onResult_inverter;
  reg        [31:0]   FpuF2iPlugin_logic_onResult_resultRaw;
  wire       [0:0]    _zz_FpuF2iPlugin_logic_onResult_expMax;
  wire       [5:0]    FpuF2iPlugin_logic_onResult_expMax;
  wire       [5:0]    FpuF2iPlugin_logic_onResult_expMin;
  wire       [31:0]   FpuF2iPlugin_logic_onResult_unsignedMin;
  reg                 FpuF2iPlugin_logic_onResult_overflow;
  wire                FpuF2iPlugin_logic_onResult_underflow;
  wire                FpuF2iPlugin_logic_onResult_isZero;
  wire                when_FpuF2iPlugin_l123;
  wire                when_FpuF2iPlugin_l136;
  wire                when_FpuF2iPlugin_l138;
  wire                when_FpuF2iPlugin_l129;
  wire       [4:0]    _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX;
  wire       [52:0]   FpuMulPlugin_logic_mulCmd_m1;
  wire       [52:0]   FpuMulPlugin_logic_mulCmd_m2;
  wire                FpuMulPlugin_logic_norm_needShift;
  reg                 FpuMulPlugin_logic_onPack_nv;
  reg        [1:0]    FpuMulPlugin_logic_onPack_mode;
  wire                when_FpuMulPlugin_l148;
  wire       [104:0]  _zz_when_AFix_l852_1;
  reg        [53:0]   _zz_FpuMulPlugin_logic_packPort_cmd_value_mantissa;
  wire                when_AFix_l852_1;
  reg                 FpuSqrtPlugin_logic_onExecute_isZero;
  wire                when_FpuSqrtPlugin_l66;
  reg                 FpuSqrtPlugin_logic_onExecute_cmdSent;
  wire                io_input_fire;
  reg                 FpuSqrtPlugin_logic_onExecute_unscheduleRequest;
  wire                FpuSqrtPlugin_logic_onExecute_freeze;
  wire       [10:0]   FpuSqrtPlugin_logic_onExecute_exp;
  wire                FpuSqrtPlugin_logic_onExecute_scrap;
  wire                FpuSqrtPlugin_logic_onExecute_negative;
  wire                when_FpuSqrtPlugin_l92;
  reg                 FpuSqrtPlugin_logic_onExecute_NV;
  wire                when_FpuSqrtPlugin_l101;
  wire                when_FpuSqrtPlugin_l105;
  wire       [0:0]    _zz_FpuXxPlugin_logic_packPort_cmd_format;
  wire                when_FpuDivPlugin_l68;
  wire                FpuDivPlugin_logic_onExecute_needShift;
  wire       [53:0]   FpuDivPlugin_logic_onExecute_mantissa;
  reg        [12:0]   _zz_FpuDivPlugin_logic_onExecute_exponent;
  wire       [12:0]   FpuDivPlugin_logic_onExecute_exponent;
  wire                FpuDivPlugin_logic_onExecute_forceOverflow;
  wire                FpuDivPlugin_logic_onExecute_infinitynan;
  wire                FpuDivPlugin_logic_onExecute_forceNan;
  wire                FpuDivPlugin_logic_onExecute_forceZero;
  wire                when_FpuDivPlugin_l102;
  wire                TrapPlugin_logic_initHold;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext_1;
  wire                when_CtrlLaneApi_l50_4;
  wire                WhiteboxerPlugin_logic_serializeds_0_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_0_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_0_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_0_microOp;
  reg                 decode_ctrls_1_up_LANE_SEL_1_regNext_1;
  wire                when_CtrlLaneApi_l50_5;
  wire                WhiteboxerPlugin_logic_serializeds_1_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_1_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_1_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_1_microOp;
  reg                 execute_ctrl0_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_6;
  wire                WhiteboxerPlugin_logic_dispatches_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_0_microOpId;
  wire                execute_lane1_ctrls_0_upIsCancel;
  wire                execute_lane1_ctrls_0_downIsCancel;
  reg                 execute_ctrl0_down_LANE_SEL_lane1_regNext;
  wire                when_CtrlLaneApi_l50_7;
  wire                WhiteboxerPlugin_logic_dispatches_1_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_1_microOpId;
  reg                 execute_ctrl2_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_8;
  wire                WhiteboxerPlugin_logic_executes_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_0_microOpId;
  reg                 execute_ctrl2_down_LANE_SEL_lane1_regNext;
  wire                when_CtrlLaneApi_l50_9;
  wire                WhiteboxerPlugin_logic_executes_1_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_1_microOpId;
  wire                WhiteboxerPlugin_logic_csr_access_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_access_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_access_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_read;
  wire                WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_access_payload_readDone;
  wire       [11:0]   BtbPlugin_logic_onForget_hash;
  wire                fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200;
  wire       [3:0]    BtbPlugin_logic_predictions;
  wire       [1:0]    BtbPlugin_logic_applyIt_chunksMask;
  wire       [1:0]    BtbPlugin_logic_applyIt_chunksTakenOh;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l233;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire                _zz_BtbPlugin_logic_applyIt_doItSlice;
  wire       [11:0]   BtbPlugin_logic_applyIt_entry_hash;
  wire       [0:0]    BtbPlugin_logic_applyIt_entry_sliceLow;
  wire       [30:0]   BtbPlugin_logic_applyIt_entry_pcTarget;
  wire                BtbPlugin_logic_applyIt_entry_isBranch;
  wire                BtbPlugin_logic_applyIt_entry_isPush;
  wire                BtbPlugin_logic_applyIt_entry_isPop;
  wire       [46:0]   _zz_BtbPlugin_logic_applyIt_entry_hash;
  reg        [30:0]   BtbPlugin_logic_applyIt_pcTarget;
  wire       [1:0]    BtbPlugin_logic_applyIt_doItSlice;
  wire                BtbPlugin_logic_applyIt_rasLogic_pushValid;
  reg        [31:0]   BtbPlugin_logic_applyIt_rasLogic_pushPc;
  wire                when_BtbPlugin_l246;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_0_history;
  wire                BtbPlugin_logic_applyIt_history_layers_0_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_1_history;
  wire                BtbPlugin_logic_applyIt_history_layers_1_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_2_history;
  wire                BtbPlugin_logic_applyIt_history_layers_2_valid;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_0_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_0_shifted;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_1_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_1_shifted;
  reg                 TrapPlugin_logic_harts_0_crsPorts_read_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_read_ready;
  reg        [1:0]    TrapPlugin_logic_harts_0_crsPorts_read_address;
  wire       [31:0]   TrapPlugin_logic_harts_0_crsPorts_read_data;
  wire                AlignerPlugin_logic_buffer_flushIt;
  wire                AlignerPlugin_logic_buffer_readers_0_firstFromBuffer;
  wire                AlignerPlugin_logic_buffer_readers_0_lastFromBuffer;
  wire       [7:0]    _zz_AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc_2;
  wire                AlignerPlugin_logic_buffer_readers_1_firstFromBuffer;
  wire                AlignerPlugin_logic_buffer_readers_1_lastFromBuffer;
  wire       [6:0]    _zz_AlignerPlugin_logic_extractors_1_ctx_instruction;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc_2;
  wire                DispatchPlugin_logic_slotsFeeds_free;
  wire                DispatchPlugin_logic_slotsFeeds_fit;
  wire                DispatchPlugin_logic_slotsFeeds_doIt;
  wire       [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid;
  wire                _zz_DispatchPlugin_logic_slots_0_ctx_valid_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid_3;
  wire       [197:0]  _zz_DispatchPlugin_logic_slots_0_ctx_valid_4;
  wire       [160:0]  _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [7:0]    _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_0;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_1;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_2;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_3;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_1;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_2;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_3;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_0_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_doIt;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_3;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_1_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_1_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_doIt;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_3;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_3;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_2_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_2_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_doIt;
  wire       [2:0]    DispatchPlugin_logic_inserter_0_oh;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane0;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane0_1;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane0_2;
  wire                DispatchPlugin_logic_inserter_0_trap;
  wire       [7:0]    _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire                when_DispatchPlugin_l439;
  wire       [3:0]    DispatchPlugin_logic_inserter_0_layerOhUnfiltred;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layer_0_0;
  wire                DispatchPlugin_logic_inserter_0_layer_0_1;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layer_1_0;
  wire                DispatchPlugin_logic_inserter_0_layer_1_1;
  wire       [1:0]    _zz_execute_ctrl0_up_lane0_LAYER_SEL_lane0;
  wire       [2:0]    DispatchPlugin_logic_inserter_1_oh;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane1;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane1_1;
  wire                _zz_execute_ctrl0_up_LANE_AGE_lane1_2;
  wire                DispatchPlugin_logic_inserter_1_trap;
  wire       [7:0]    _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire                when_DispatchPlugin_l439_1;
  wire       [3:0]    DispatchPlugin_logic_inserter_1_layerOhUnfiltred;
  wire       [0:0]    DispatchPlugin_logic_inserter_1_layer_0_0;
  wire                DispatchPlugin_logic_inserter_1_layer_0_1;
  wire       [0:0]    DispatchPlugin_logic_inserter_1_layer_1_0;
  wire                DispatchPlugin_logic_inserter_1_layer_1_1;
  wire       [1:0]    _zz_execute_ctrl0_up_lane1_LAYER_SEL_lane1;
  wire                decode_logic_flushes_0_onLanes_0_doIt;
  wire                decode_logic_flushes_0_onLanes_1_doIt;
  wire                decode_logic_flushes_1_onLanes_0_doIt;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt;
  wire                decode_logic_flushes_1_onLanes_1_doIt;
  wire                execute_lane1_bypasser_integer_RS1_port_valid;
  wire       [4:0]    execute_lane1_bypasser_integer_RS1_port_address;
  wire       [31:0]   execute_lane1_bypasser_integer_RS1_port_data;
  reg                 TrapPlugin_logic_harts_0_crsPorts_write_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_write_ready;
  reg        [1:0]    TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [31:0]   TrapPlugin_logic_harts_0_crsPorts_write_data;
  reg                 TrapPlugin_logic_harts_0_interrupt_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
  wire                when_TrapPlugin_l201;
  wire                when_TrapPlugin_l207;
  wire                when_TrapPlugin_l207_1;
  wire                when_TrapPlugin_l207_2;
  reg                 TrapPlugin_logic_harts_0_interrupt_validBuffer;
  wire                TrapPlugin_logic_harts_0_interrupt_pendingInterrupt;
  wire                when_TrapPlugin_l226;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
  wire       [38:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  reg                 TrapPlugin_logic_harts_0_trap_pending_state_exception;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_state_tval;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_pending_state_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_state_arg;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_pc;
  reg        [11:0]   TrapPlugin_logic_harts_0_trap_pending_history;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_exception_code;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_exception_targetPrivilege;
  wire                execute_lane1_ctrls_5_upIsCancel;
  wire                execute_lane1_ctrls_5_downIsCancel;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_trigger_oh;
  wire                TrapPlugin_logic_harts_0_trap_trigger_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_pc;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_pc_1;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_trap;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_whitebox_code;
  reg                 TrapPlugin_logic_harts_0_trap_historyPort_valid;
  wire       [11:0]   TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  reg                 TrapPlugin_logic_harts_0_trap_pcPort_valid;
  wire                TrapPlugin_logic_harts_0_trap_pcPort_payload_fault;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantExit;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wantStart;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantKill;
  wire                TrapPlugin_logic_harts_0_trap_fsm_inflightTrap;
  wire                TrapPlugin_logic_harts_0_trap_fsm_holdPort;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wfi;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege;
  wire                TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
  wire                TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_jumpOffset;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug;
  wire                TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg;
  wire                when_TrapPlugin_l556;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_readed;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege;
  wire                PcPlugin_logic_forcedSpawn;
  reg        [9:0]    PcPlugin_logic_harts_0_self_id;
  wire                PcPlugin_logic_harts_0_self_flow_valid;
  wire                PcPlugin_logic_harts_0_self_flow_payload_fault;
  wire       [31:0]   PcPlugin_logic_harts_0_self_flow_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid;
  reg                 PcPlugin_logic_harts_0_self_increment;
  reg                 PcPlugin_logic_harts_0_self_fault;
  reg        [31:0]   PcPlugin_logic_harts_0_self_state;
  wire       [31:0]   PcPlugin_logic_harts_0_self_pc;
  wire                PcPlugin_logic_harts_0_aggregator_valids_0;
  wire                PcPlugin_logic_harts_0_aggregator_valids_1;
  wire                PcPlugin_logic_harts_0_aggregator_valids_2;
  wire                PcPlugin_logic_harts_0_aggregator_valids_3;
  wire                PcPlugin_logic_harts_0_aggregator_valids_4;
  wire                PcPlugin_logic_harts_0_aggregator_valids_5;
  wire                PcPlugin_logic_harts_0_aggregator_valids_6;
  wire       [6:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_3;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_5;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_6;
  reg        [6:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh_7;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_8;
  wire       [6:0]    PcPlugin_logic_harts_0_aggregator_oh;
  (* keep , syn_keep *) wire       [31:0]   PcPlugin_logic_harts_0_aggregator_target /* synthesis syn_keep = 1 */ ;
  wire                PcPlugin_logic_harts_0_aggregator_fault;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_3;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_4;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_5;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_fault_1;
  wire                when_PcPlugin_l80;
  wire                PcPlugin_logic_harts_0_holdComb;
  reg                 PcPlugin_logic_harts_0_holdReg;
  wire                PcPlugin_logic_harts_0_output_valid;
  wire                PcPlugin_logic_harts_0_output_ready;
  reg        [31:0]   PcPlugin_logic_harts_0_output_payload_pc;
  wire                PcPlugin_logic_harts_0_output_payload_fault;
  wire                PcPlugin_logic_harts_0_output_fire;
  wire                PcPlugin_logic_holdHalter_doIt;
  wire                fetch_logic_ctrls_0_haltRequest_PcPlugin_l133;
  wire                CsrAccessPlugin_logic_fsm_wantExit;
  reg                 CsrAccessPlugin_logic_fsm_wantStart;
  wire                CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_2047;
  reg                 REG_CSR_1952;
  reg                 REG_CSR_1953;
  reg                 REG_CSR_1954;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_768;
  reg                 REG_CSR_834;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_3;
  reg                 REG_CSR_2;
  reg                 REG_CSR_1;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  reg                 REG_CSR_FpuCsrPlugin_logic_csrDirty;
  reg                 REG_CSR_CsrRamPlugin_csrMapper_selFilter;
  reg                 REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  reg                 CsrAccessPlugin_logic_fsm_interface_read;
  reg                 CsrAccessPlugin_logic_fsm_interface_write;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_interface_rs1;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_aluInput;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_csrValue;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  wire       [15:0]   CsrAccessPlugin_logic_fsm_interface_uopId;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_interface_uop;
  wire                CsrAccessPlugin_logic_fsm_interface_doImm;
  wire                CsrAccessPlugin_logic_fsm_interface_doMask;
  wire                CsrAccessPlugin_logic_fsm_interface_doClear;
  wire       [4:0]    CsrAccessPlugin_logic_fsm_interface_rdPhys;
  wire                CsrAccessPlugin_logic_fsm_interface_rdEnable;
  reg                 CsrAccessPlugin_logic_fsm_interface_fire;
  wire       [11:0]   CsrAccessPlugin_logic_fsm_inject_csrAddress;
  wire                CsrAccessPlugin_logic_fsm_inject_immZero;
  wire                CsrAccessPlugin_logic_fsm_inject_srcZero;
  wire                CsrAccessPlugin_logic_fsm_inject_csrWrite;
  wire                CsrAccessPlugin_logic_fsm_inject_csrRead;
  wire                COMB_CSR_2047;
  wire                COMB_CSR_1952;
  wire                COMB_CSR_1953;
  wire                COMB_CSR_1954;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_768;
  wire                COMB_CSR_834;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_3;
  wire                COMB_CSR_2;
  wire                COMB_CSR_1;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  wire                COMB_CSR_FpuCsrPlugin_logic_csrDirty;
  wire                COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  wire                CsrAccessPlugin_logic_fsm_inject_implemented;
  wire                CsrAccessPlugin_logic_fsm_inject_onDecodeDo;
  wire                when_CsrAccessPlugin_l155;
  wire                CsrAccessPlugin_logic_fsm_inject_trap;
  reg                 CsrAccessPlugin_logic_fsm_inject_unfreeze;
  wire                CsrAccessPlugin_logic_fsm_inject_freeze;
  reg                 CsrAccessPlugin_logic_fsm_inject_flushReg;
  wire                when_CsrAccessPlugin_l197;
  reg                 CsrAccessPlugin_logic_fsm_inject_sampled;
  reg                 CsrAccessPlugin_logic_fsm_inject_trapReg;
  reg                 CsrAccessPlugin_logic_fsm_inject_busTrapReg;
  reg        [3:0]    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  wire                when_CsrAccessPlugin_l252;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l346;
  wire                when_CsrAccessPlugin_l346_1;
  wire                when_CsrAccessPlugin_l346_2;
  wire                when_CsrAccessPlugin_l346_3;
  wire                when_CsrAccessPlugin_l346_4;
  wire       [4:0]    _zz_FpuCsrPlugin_api_flags_NX;
  wire                when_CsrAccessPlugin_l346_5;
  wire                when_CsrAccessPlugin_l346_6;
  wire       [4:0]    _zz_FpuCsrPlugin_api_flags_NX_1;
  wire                when_CsrAccessPlugin_l343;
  wire                when_CsrAccessPlugin_l343_1;
  wire                when_CsrAccessPlugin_l346_7;
  wire                when_CsrAccessPlugin_l343_2;
  reg        [11:0]   HistoryPlugin_logic_onFetch_value;
  reg        [11:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire                HistoryPlugin_logic_onFetch_ports_0_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_0_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_1_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire       [0:0]    HistoryPlugin_logic_onFetch_ports_1_payload_age;
  wire       [12:0]   _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_2_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_2_payload_history;
  wire       [0:0]    HistoryPlugin_logic_onFetch_ports_2_payload_age;
  wire       [12:0]   _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_3_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_3_payload_history;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [1:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [31:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire                _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  wire                _zz_CsrRamPlugin_csrMapper_write_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel;
  wire       [0:0]    CsrRamPlugin_logic_readLogic_sel;
  wire                CsrRamPlugin_logic_readLogic_port_cmd_valid;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [31:0]   CsrRamPlugin_logic_readLogic_port_rsp;
  reg        [1:0]    CsrRamPlugin_logic_readLogic_ohReg;
  reg                 CsrRamPlugin_logic_readLogic_busy;
  reg        [2:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                execute_lane0_bypasser_integer_RS1_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS1_port_address;
  wire       [31:0]   execute_lane0_bypasser_integer_RS1_port_data;
  reg        [8:0]    execute_lane0_bypasser_integer_RS1_bypassEnables;
  wire       [8:0]    _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8;
  reg        [8:0]    _zz_execute_lane0_bypasser_integer_RS1_sel;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7;
  wire       [8:0]    execute_lane0_bypasser_integer_RS1_sel;
  wire       [7:0]    _zz_execute_ctrl1_down_integer_RS1_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS1_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit;
  wire       [2:0]    execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits;
  wire       [3:0]    _zz_execute_ctrl2_integer_RS1_lane0_bypass;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit;
  wire                execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit;
  wire       [1:0]    execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits;
  wire       [2:0]    _zz_execute_ctrl3_integer_RS1_lane0_bypass;
  wire                execute_lane0_bypasser_integer_RS2_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS2_port_address;
  wire       [31:0]   execute_lane0_bypasser_integer_RS2_port_data;
  reg        [8:0]    execute_lane0_bypasser_integer_RS2_bypassEnables;
  wire       [8:0]    _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8;
  reg        [8:0]    _zz_execute_lane0_bypasser_integer_RS2_sel;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7;
  wire       [8:0]    execute_lane0_bypasser_integer_RS2_sel;
  wire       [7:0]    _zz_execute_ctrl1_down_integer_RS2_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS2_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196_1;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit;
  wire       [2:0]    execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits;
  wire       [3:0]    _zz_execute_ctrl2_integer_RS2_lane0_bypass;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit;
  wire                execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit;
  wire       [1:0]    execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits;
  wire       [2:0]    _zz_execute_ctrl3_integer_RS2_lane0_bypass;
  wire                execute_lane0_bypasser_float_RS1_port_valid;
  wire       [4:0]    execute_lane0_bypasser_float_RS1_port_address;
  wire       [63:0]   execute_lane0_bypasser_float_RS1_port_data;
  reg        [9:0]    execute_lane0_bypasser_float_RS1_bypassEnables;
  wire                execute_lane0_ctrls_12_upIsCancel;
  wire                execute_lane0_ctrls_12_downIsCancel;
  wire       [9:0]    _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_4;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_5;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_6;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_7;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_8;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_bools_9;
  reg        [9:0]    _zz_execute_lane0_bypasser_float_RS1_sel;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_5;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_6;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_7;
  wire                execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_7;
  wire       [9:0]    execute_lane0_bypasser_float_RS1_sel;
  wire                execute_lane0_bypasser_float_RS2_port_valid;
  wire       [4:0]    execute_lane0_bypasser_float_RS2_port_address;
  wire       [63:0]   execute_lane0_bypasser_float_RS2_port_data;
  reg        [9:0]    execute_lane0_bypasser_float_RS2_bypassEnables;
  wire       [9:0]    _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_4;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_5;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_6;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_7;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_8;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_bools_9;
  reg        [9:0]    _zz_execute_lane0_bypasser_float_RS2_sel;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_5;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_6;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_7;
  wire                execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_7;
  wire       [9:0]    execute_lane0_bypasser_float_RS2_sel;
  wire                execute_lane0_bypasser_float_RS3_port_valid;
  wire       [4:0]    execute_lane0_bypasser_float_RS3_port_address;
  wire       [63:0]   execute_lane0_bypasser_float_RS3_port_data;
  reg        [9:0]    execute_lane0_bypasser_float_RS3_bypassEnables;
  wire       [9:0]    _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_4;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_5;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_6;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_7;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_8;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_bools_9;
  reg        [9:0]    _zz_execute_lane0_bypasser_float_RS3_sel;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_5;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_6;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_7;
  wire                execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_7;
  wire       [9:0]    execute_lane0_bypasser_float_RS3_sel;
  wire                execute_lane0_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_2_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_3_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_3_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_3_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_3_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_4_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_4_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_4_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_4_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_5_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_5_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_5_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_5_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_6_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_6_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_6_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_6_port_payload_commit;
  wire       [32:0]   execute_lane0_logic_decoding_decodingBits;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_4;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_5;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_6;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_7;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_8;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_9;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_11;
  wire                _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_12;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_13;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_14;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_15;
  wire                _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                _zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire                _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire                _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0;
  wire                _zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1;
  wire                _zz_execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_1;
  wire                _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  wire                _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0;
  wire                _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [1:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire       [1:0]    _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3;
  wire                when_ExecuteLanePlugin_l306;
  wire                when_ExecuteLanePlugin_l306_1;
  wire                when_ExecuteLanePlugin_l306_2;
  wire                when_ExecuteLanePlugin_l306_3;
  wire                when_ExecuteLanePlugin_l306_4;
  wire                when_FpuFlagsWritebackPlugin_l96;
  wire                WhiteboxerPlugin_logic_csr_port_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_port_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_port_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_read;
  wire                WhiteboxerPlugin_logic_csr_port_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_port_payload_readDone;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_3_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_3_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_4_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_4_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_5_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_5_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_6_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_6_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_6_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_7_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_7_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_7_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_8_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_8_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_8_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_9_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_9_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_9_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_10_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_10_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_10_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_11_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_11_payload_uopId;
  wire       [63:0]   WhiteboxerPlugin_logic_rfWrites_ports_11_payload_data;
  wire                WhiteboxerPlugin_logic_completions_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_0_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_4_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_4_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_4_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_5_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_5_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_5_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_6_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_6_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_6_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_6_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_7_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_7_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_7_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_7_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_8_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_8_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_8_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_8_payload_commit;
  wire                fetch_logic_flushes_0_doIt;
  wire                fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48;
  wire                fetch_logic_flushes_1_doIt;
  wire                fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50;
  reg        [8:0]    execute_lane1_bypasser_integer_RS1_bypassEnables;
  wire       [8:0]    _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8;
  reg        [8:0]    _zz_execute_lane1_bypasser_integer_RS1_sel;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6;
  wire                execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7;
  wire       [8:0]    execute_lane1_bypasser_integer_RS1_sel;
  wire       [7:0]    _zz_execute_ctrl1_down_integer_RS1_lane1;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS1_lane1_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196_2;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit;
  wire       [2:0]    execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits;
  wire       [3:0]    _zz_execute_ctrl2_integer_RS1_lane1_bypass;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit;
  wire                execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit;
  wire       [1:0]    execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits;
  wire       [2:0]    _zz_execute_ctrl3_integer_RS1_lane1_bypass;
  wire                execute_lane1_bypasser_integer_RS2_port_valid;
  wire       [4:0]    execute_lane1_bypasser_integer_RS2_port_address;
  wire       [31:0]   execute_lane1_bypasser_integer_RS2_port_data;
  reg        [8:0]    execute_lane1_bypasser_integer_RS2_bypassEnables;
  wire       [8:0]    _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8;
  reg        [8:0]    _zz_execute_lane1_bypasser_integer_RS2_sel;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6;
  wire                execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7;
  wire       [8:0]    execute_lane1_bypasser_integer_RS2_sel;
  wire       [7:0]    _zz_execute_ctrl1_down_integer_RS2_lane1;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS2_lane1_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196_3;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit;
  wire       [2:0]    execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits;
  wire       [3:0]    _zz_execute_ctrl2_integer_RS2_lane1_bypass;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit;
  wire                execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit;
  wire       [1:0]    execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits;
  wire       [2:0]    _zz_execute_ctrl3_integer_RS2_lane1_bypass;
  wire                execute_lane1_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane1_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane1_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane1_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane1_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane1_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane1_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane1_logic_completions_onCtrl_1_port_payload_commit;
  wire       [32:0]   execute_lane1_logic_decoding_decodingBits;
  wire                _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
  wire                _zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1;
  wire                _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire                _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
  wire                _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  wire       [1:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire       [1:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  wire       [1:0]    _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  wire                _zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2;
  wire       [1:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  wire       [1:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3;
  wire       [1:0]    _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4;
  wire                when_ExecuteLanePlugin_l306_5;
  wire                when_ExecuteLanePlugin_l306_6;
  wire                when_ExecuteLanePlugin_l306_7;
  wire                when_ExecuteLanePlugin_l306_8;
  wire                when_ExecuteLanePlugin_l306_9;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_uopId;
  reg        [5:0]    integer_RegFilePlugin_logic_initalizer_counter;
  wire                integer_RegFilePlugin_logic_initalizer_done;
  wire                when_RegFilePlugin_l132;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [4:0]    integer_write_0_address /* verilator public */ ;
  wire       [31:0]   integer_write_0_data /* verilator public */ ;
  wire       [15:0]   integer_write_0_uopId /* verilator public */ ;
  wire                integer_write_1_valid /* verilator public */ ;
  wire       [4:0]    integer_write_1_address /* verilator public */ ;
  wire       [31:0]   integer_write_1_data /* verilator public */ ;
  wire       [15:0]   integer_write_1_uopId /* verilator public */ ;
  wire                float_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [4:0]    float_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [63:0]   float_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [15:0]   float_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  reg        [5:0]    float_RegFilePlugin_logic_initalizer_counter;
  wire                float_RegFilePlugin_logic_initalizer_done;
  wire                when_RegFilePlugin_l132_1;
  wire                float_write_0_valid /* verilator public */ ;
  wire       [4:0]    float_write_0_address /* verilator public */ ;
  wire       [63:0]   float_write_0_data /* verilator public */ ;
  wire       [15:0]   float_write_0_uopId /* verilator public */ ;
  wire                WhiteboxerPlugin_logic_completions_ports_9_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_9_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_9_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_9_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_10_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_10_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_10_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_10_payload_commit;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_1;
  wire                WhiteboxerPlugin_logic_commits_ports_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_uop;
  wire                WhiteboxerPlugin_logic_commits_ports_1_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_1_oh_1;
  wire                WhiteboxerPlugin_logic_commits_ports_1_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_1_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_1_uop;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_valid;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_1_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_2_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_3_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_4_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_5_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_6_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_6_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_6_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_6_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_7_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_7_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_7_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_7_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_8_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_8_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_8_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_8_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_9_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_9_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_9_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_9_payload_self;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  wire       [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  wire       [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_pcOnLastSlice;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                WhiteboxerPlugin_logic_loadExecute_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_loadExecute_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_loadExecute_size;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_address;
  reg        [63:0]   WhiteboxerPlugin_logic_loadExecute_data;
  wire                WhiteboxerPlugin_logic_storeCommit_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeCommit_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_storeCommit_storeId;
  wire       [1:0]    WhiteboxerPlugin_logic_storeCommit_size;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_address;
  wire       [63:0]   WhiteboxerPlugin_logic_storeCommit_data;
  wire                WhiteboxerPlugin_logic_storeCommit_amo;
  wire                WhiteboxerPlugin_logic_storeConditional_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeConditional_uopId;
  wire                WhiteboxerPlugin_logic_storeConditional_miss;
  wire                WhiteboxerPlugin_logic_storeBroadcast_fire;
  wire       [11:0]   WhiteboxerPlugin_logic_storeBroadcast_storeId;
  wire       [0:0]    WhiteboxerPlugin_logic_wfi;
  wire                WhiteboxerPlugin_logic_perf_executeFreezed;
  wire                WhiteboxerPlugin_logic_perf_dispatchHazards;
  wire       [1:0]    WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [1:0]    WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  reg                 _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  wire                when_Utils_l593;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  wire                when_Utils_l593_1;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  wire                when_Utils_l593_2;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  wire                when_Utils_l593_3;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  wire                when_Utils_l593_4;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  wire                when_Utils_l593_5;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  wire                when_Utils_l593_6;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  wire                WhiteboxerPlugin_logic_trap_ports_0_valid;
  wire                WhiteboxerPlugin_logic_trap_ports_0_interrupt;
  wire       [3:0]    WhiteboxerPlugin_logic_trap_ports_0_cause;
  wire                fetch_logic_ctrls_2_up_forgetOne;
  wire                fetch_logic_ctrls_1_up_forgetOne;
  wire                when_CtrlLink_l191;
  wire                when_CtrlLink_l198;
  wire                when_StageLink_l71_3;
  wire                when_DecodePipelinePlugin_l70;
  wire                when_DecodePipelinePlugin_l70_1;
  reg        [1:0]    LsuPlugin_logic_flusher_stateReg;
  reg        [1:0]    LsuPlugin_logic_flusher_stateNext;
  wire                when_LsuPlugin_l363;
  wire                when_LsuPlugin_l371;
  wire                LsuPlugin_logic_flusher_onExit_IDLE;
  wire                LsuPlugin_logic_flusher_onExit_SB_DRAIN;
  wire                LsuPlugin_logic_flusher_onExit_CMD;
  wire                LsuPlugin_logic_flusher_onExit_COMPLETION;
  wire                LsuPlugin_logic_flusher_onEntry_IDLE;
  wire                LsuPlugin_logic_flusher_onEntry_SB_DRAIN;
  wire                LsuPlugin_logic_flusher_onEntry_CMD;
  wire                LsuPlugin_logic_flusher_onEntry_COMPLETION;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateReg;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateNext;
  wire                when_TrapPlugin_l409;
  wire                when_TrapPlugin_l654;
  wire       [1:0]    switch_TrapPlugin_l655;
  wire                when_TrapPlugin_l362;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_COMPUTE;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_COMPUTE;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateReg;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateNext;
  wire                when_CsrAccessPlugin_l296;
  wire                when_CsrAccessPlugin_l325;
  wire                when_CsrAccessPlugin_l212;
  wire                CsrAccessPlugin_logic_fsm_onExit_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onExit_READ;
  wire                CsrAccessPlugin_logic_fsm_onExit_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onExit_COMPLETION;
  wire                CsrAccessPlugin_logic_fsm_onEntry_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_READ;
  wire                CsrAccessPlugin_logic_fsm_onEntry_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_COMPLETION;
  `ifndef SYNTHESIS
  reg [47:0] execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [47:0] execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [23:0] execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string;
  reg [191:0] execute_ctrl4_down_FpuUtils_FORMAT_lane0_string;
  reg [47:0] execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [47:0] execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [47:0] execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [23:0] execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string;
  reg [191:0] execute_ctrl5_up_FpuUtils_FORMAT_lane0_string;
  reg [47:0] execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [39:0] execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [47:0] execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [47:0] execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [47:0] execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [23:0] execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string;
  reg [39:0] execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [191:0] execute_ctrl4_up_FpuUtils_FORMAT_lane0_string;
  reg [31:0] execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [47:0] execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [47:0] execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [47:0] execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [23:0] execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string;
  reg [39:0] execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [55:0] execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [191:0] execute_ctrl3_up_FpuUtils_FORMAT_lane0_string;
  reg [31:0] execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string;
  reg [55:0] execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [191:0] execute_ctrl2_up_FpuUtils_FORMAT_lane0_string;
  reg [31:0] execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string;
  reg [55:0] execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [191:0] execute_ctrl1_down_FpuUtils_FORMAT_lane0_string;
  reg [31:0] execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [47:0] execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [23:0] execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string;
  reg [191:0] execute_ctrl5_down_FpuUtils_FORMAT_lane0_string;
  reg [47:0] execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [47:0] execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [47:0] execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [23:0] execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string;
  reg [47:0] execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [55:0] execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [55:0] execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [47:0] execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [191:0] execute_ctrl3_down_FpuUtils_FORMAT_lane0_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string;
  reg [47:0] execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string;
  reg [191:0] execute_ctrl2_down_FpuUtils_FORMAT_lane0_string;
  reg [31:0] execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [23:0] FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string;
  reg [47:0] FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string;
  reg [191:0] FpuPackerPlugin_logic_pip_node_2_s0_FORMAT_string;
  reg [23:0] FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string;
  reg [191:0] FpuPackerPlugin_logic_pip_node_1_s0_FORMAT_string;
  reg [47:0] FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string;
  reg [23:0] FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string;
  reg [191:0] FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string;
  reg [47:0] FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string;
  reg [23:0] execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string;
  reg [31:0] execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [23:0] FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string;
  reg [191:0] FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT_string;
  reg [23:0] FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string;
  reg [191:0] FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT_string;
  reg [23:0] FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string;
  reg [191:0] FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT_string;
  reg [23:0] FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string;
  reg [191:0] FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string;
  reg [23:0] FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string;
  reg [191:0] FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string;
  reg [79:0] execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string;
  reg [39:0] execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [47:0] FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuUnpackerPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuAddPlugin_logic_addPort_cmd_rs1_mode_string;
  reg [47:0] FpuAddPlugin_logic_addPort_cmd_rs2_mode_string;
  reg [191:0] FpuAddPlugin_logic_addPort_cmd_format_string;
  reg [23:0] FpuAddPlugin_logic_addPort_cmd_roundMode_string;
  reg [47:0] FpuMulPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuMulPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuMulPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuSqrtPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuSqrtPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuSqrtPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuXxPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuXxPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuXxPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuDivPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuDivPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuDivPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuMulPlugin_logic_addPort_cmd_rs1_mode_string;
  reg [47:0] FpuMulPlugin_logic_addPort_cmd_rs2_mode_string;
  reg [191:0] FpuMulPlugin_logic_addPort_cmd_format_string;
  reg [23:0] FpuMulPlugin_logic_addPort_cmd_roundMode_string;
  reg [47:0] FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string;
  reg [191:0] FpuAddSharedPlugin_logic_packPort_cmd_format_string;
  reg [23:0] FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string;
  reg [47:0] FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string;
  reg [47:0] FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string;
  reg [47:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string;
  reg [47:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string;
  reg [47:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string;
  reg [47:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string;
  reg [191:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string;
  reg [191:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1_string;
  reg [23:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string;
  reg [23:0] _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string;
  reg [23:0] _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string;
  reg [95:0] LsuPlugin_logic_onAddress0_ls_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_flush_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_sb_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_0_mode_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_1_mode_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_2_mode_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_3_mode_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_4_mode_string;
  reg [47:0] FpuPackerPlugin_logic_s0_remapped_5_mode_string;
  reg [47:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string;
  reg [47:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string;
  reg [191:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string;
  reg [191:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_string;
  reg [23:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string;
  reg [23:0] _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string;
  reg [47:0] _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string;
  reg [47:0] FpuMulPlugin_logic_onPack_mode_string;
  reg [191:0] _zz_FpuXxPlugin_logic_packPort_cmd_format_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string;
  reg [191:0] _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_string;
  reg [191:0] _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_string;
  reg [191:0] _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2_string;
  reg [55:0] _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string;
  reg [55:0] _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1_string;
  reg [55:0] _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string;
  reg [39:0] _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [39:0] _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string;
  reg [39:0] _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string;
  reg [39:0] _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string;
  reg [39:0] _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string;
  reg [39:0] _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string;
  reg [39:0] _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string;
  reg [79:0] LsuPlugin_logic_flusher_stateReg_string;
  reg [79:0] LsuPlugin_logic_flusher_stateNext_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateReg_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateNext_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateNext_string;
  `endif

  (* ram_style = "distributed" *) reg [30:0] BtbPlugin_logic_ras_mem_stack [0:3];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol0 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol1 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol2 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol3 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol4 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol5 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol6 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol7 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol8 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol9 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol10 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol11 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol12 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol13 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol14 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol15 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol16 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol17 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol18 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol19 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol20 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol21 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol22 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol23 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol24 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol25 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol26 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol27 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol28 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol29 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol30 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol31 [0:127];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_8;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_9;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_10;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_11;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_12;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_13;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_14;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_15;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_16;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_17;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_18;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_19;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_20;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_21;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_22;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_23;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_24;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_25;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_26;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_27;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_28;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_29;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_30;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_31;
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol0 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol1 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol2 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol3 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol4 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol5 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol6 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol7 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol8 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol9 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol10 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol11 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol12 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol13 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol14 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol15 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol16 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol17 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol18 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol19 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol20 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol21 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol22 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol23 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol24 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol25 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol26 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol27 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol28 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol29 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol30 [0:127];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol31 [0:127];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_8;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_9;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_10;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_11;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_12;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_13;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_14;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_15;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_16;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_17;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_18;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_19;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_20;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_21;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_22;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_23;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_24;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_25;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_26;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_27;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_28;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_29;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_30;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_31;
  reg [21:0] LsuL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_1_mem [0:63];
  reg [2:0] LsuL1Plugin_logic_shared_mem [0:63];
  reg [255:0] LsuL1Plugin_logic_writeback_victimBuffer [0:3];
  reg [51:0] PrefetcherRptPlugin_logic_storage_ram [0:127];
  reg [255:0] FetchL1Plugin_logic_banks_0_mem [0:127];
  reg [255:0] FetchL1Plugin_logic_banks_1_mem [0:127];
  reg [21:0] FetchL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_1_mem [0:63];
  reg [0:0] FetchL1Plugin_logic_plru_mem [0:63];
  reg [7:0] GSharePlugin_logic_mem_banks_0 [0:3];
  (* ram_style = "block" *) reg [46:0] BtbPlugin_logic_mem_symbol0 [0:127];
  (* ram_style = "block" *) reg [46:0] BtbPlugin_logic_mem_symbol1 [0:127];
  reg [46:0] _zz_BtbPlugin_logic_memsymbol_read;
  reg [46:0] _zz_BtbPlugin_logic_memsymbol_read_1;
  reg [109:0] LsuPlugin_logic_storeBuffer_ops_mem [0:31];
  reg [31:0] CsrRamPlugin_logic_mem [0:3];
  function [1:0] zz_FetchL1Plugin_logic_trapPort_payload_arg(input dummy);
    begin
      zz_FetchL1Plugin_logic_trapPort_payload_arg = 2'b00;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[1 : 0] = 2'b10;
    end
  endfunction
  wire [1:0] _zz_71;

  assign _zz_when = _zz_when_1[1];
  assign _zz_when_3 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[0];
  assign _zz_when_4 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[1];
  assign _zz_when_5 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[2];
  assign _zz_when_6 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[3];
  assign _zz_when_7 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[4];
  assign _zz_when_8 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[5];
  assign _zz_when_9 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[6];
  assign _zz_when_10 = LsuPlugin_logic_storeBuffer_push_payload_slotOh[7];
  assign _zz_early0_IntAluPlugin_logic_alu_result = (early0_IntAluPlugin_logic_alu_bitwise | _zz_early0_IntAluPlugin_logic_alu_result_1);
  assign _zz_early0_IntAluPlugin_logic_alu_result_1 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_2 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_early0_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_3 = _zz_early0_IntAluPlugin_logic_alu_result_4;
  assign _zz_early0_IntAluPlugin_logic_alu_result_5 = execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  assign _zz_early0_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_early0_IntAluPlugin_logic_alu_result_5};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[4 : 0];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[0],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[1],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[2],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[3],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[4],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[5],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[6],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[7],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[8],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early0_BarrelShifterPlugin_logic_shift_shifted_1) >>> early0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 && execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]),early0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched = {early0_BarrelShifterPlugin_logic_shift_shifted[0],{early0_BarrelShifterPlugin_logic_shift_shifted[1],{early0_BarrelShifterPlugin_logic_shift_shifted[2],{early0_BarrelShifterPlugin_logic_shift_shifted[3],{early0_BarrelShifterPlugin_logic_shift_shifted[4],{early0_BarrelShifterPlugin_logic_shift_shifted[5],{early0_BarrelShifterPlugin_logic_shift_shifted[6],{early0_BarrelShifterPlugin_logic_shift_shifted[7],{early0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_2,_zz_early0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[0 : 0];
  assign _zz_LsuL1Plugin_logic_refill_free_1 = (_zz_LsuL1Plugin_logic_refill_free & (~ _zz_LsuL1Plugin_logic_refill_free_2));
  assign _zz_LsuL1Plugin_logic_refill_free_2 = (_zz_LsuL1Plugin_logic_refill_free - 2'b01);
  assign _zz_LsuL1Plugin_logic_writeback_free_1 = (_zz_LsuL1Plugin_logic_writeback_free & (~ _zz_LsuL1Plugin_logic_writeback_free_2));
  assign _zz_LsuL1Plugin_logic_writeback_free_2 = (_zz_LsuL1Plugin_logic_writeback_free - 2'b01);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite = ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault)) : 1'b0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault)) : 1'b0));
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty = (2'b01 <<< LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[0 : 0];
  assign _zz_PrefetcherRptPlugin_logic_counter = (PrefetcherRptPlugin_logic_counter + _zz_PrefetcherRptPlugin_logic_counter_1);
  assign _zz_PrefetcherRptPlugin_logic_counter_2 = PrefetcherRptPlugin_logic_pip2_node_0_isFiring;
  assign _zz_PrefetcherRptPlugin_logic_counter_1 = {2'd0, _zz_PrefetcherRptPlugin_logic_counter_2};
  assign _zz_PrefetcherRptPlugin_logic_pip2_node_0_MUL = {1'b0,PrefetcherRptPlugin_logic_advanceAt};
  assign _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR = ($signed(_zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_1) + $signed(_zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_2));
  assign _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_1 = PrefetcherRptPlugin_logic_pip2_node_1_CMD_address;
  assign _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR_2 = {{16{PrefetcherRptPlugin_logic_pip2_node_1_MUL[15]}}, PrefetcherRptPlugin_logic_pip2_node_1_MUL};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = {31'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = {31'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1};
  assign _zz_late0_IntAluPlugin_logic_alu_result = (late0_IntAluPlugin_logic_alu_bitwise | _zz_late0_IntAluPlugin_logic_alu_result_1);
  assign _zz_late0_IntAluPlugin_logic_alu_result_1 = (execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 ? execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 : 32'h0);
  assign _zz_late0_IntAluPlugin_logic_alu_result_2 = (execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_late0_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_late0_IntAluPlugin_logic_alu_result_3 = _zz_late0_IntAluPlugin_logic_alu_result_4;
  assign _zz_late0_IntAluPlugin_logic_alu_result_5 = execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
  assign _zz_late0_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_late0_IntAluPlugin_logic_alu_result_5};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[4 : 0];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[0],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[1],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[2],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[3],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[4],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[5],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[6],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[7],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[8],{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_late0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_late0_BarrelShifterPlugin_logic_shift_shifted_1) >>> late0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_late0_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0 && execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]),late0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched = {late0_BarrelShifterPlugin_logic_shift_shifted[0],{late0_BarrelShifterPlugin_logic_shift_shifted[1],{late0_BarrelShifterPlugin_logic_shift_shifted[2],{late0_BarrelShifterPlugin_logic_shift_shifted[3],{late0_BarrelShifterPlugin_logic_shift_shifted[4],{late0_BarrelShifterPlugin_logic_shift_shifted[5],{late0_BarrelShifterPlugin_logic_shift_shifted[6],{late0_BarrelShifterPlugin_logic_shift_shifted[7],{late0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_late0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_late0_BarrelShifterPlugin_logic_shift_patched_2,_zz_late0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_early1_IntAluPlugin_logic_alu_result = (early1_IntAluPlugin_logic_alu_bitwise | _zz_early1_IntAluPlugin_logic_alu_result_1);
  assign _zz_early1_IntAluPlugin_logic_alu_result_1 = (execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 ? execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 : 32'h0);
  assign _zz_early1_IntAluPlugin_logic_alu_result_2 = (execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1 ? _zz_early1_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_early1_IntAluPlugin_logic_alu_result_3 = _zz_early1_IntAluPlugin_logic_alu_result_4;
  assign _zz_early1_IntAluPlugin_logic_alu_result_5 = execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
  assign _zz_early1_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_early1_IntAluPlugin_logic_alu_result_5};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[4 : 0];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[0],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[1],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[2],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[3],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[4],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[5],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[6],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[7],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[8],{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early1_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early1_BarrelShifterPlugin_logic_shift_shifted_1) >>> early1_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early1_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1 && execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]),early1_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched = {early1_BarrelShifterPlugin_logic_shift_shifted[0],{early1_BarrelShifterPlugin_logic_shift_shifted[1],{early1_BarrelShifterPlugin_logic_shift_shifted[2],{early1_BarrelShifterPlugin_logic_shift_shifted[3],{early1_BarrelShifterPlugin_logic_shift_shifted[4],{early1_BarrelShifterPlugin_logic_shift_shifted[5],{early1_BarrelShifterPlugin_logic_shift_shifted[6],{early1_BarrelShifterPlugin_logic_shift_shifted[7],{early1_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early1_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early1_BarrelShifterPlugin_logic_shift_patched_2,_zz_early1_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_late1_IntAluPlugin_logic_alu_result = (late1_IntAluPlugin_logic_alu_bitwise | _zz_late1_IntAluPlugin_logic_alu_result_1);
  assign _zz_late1_IntAluPlugin_logic_alu_result_1 = (execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 ? execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 : 32'h0);
  assign _zz_late1_IntAluPlugin_logic_alu_result_2 = (execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1 ? _zz_late1_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_late1_IntAluPlugin_logic_alu_result_3 = _zz_late1_IntAluPlugin_logic_alu_result_4;
  assign _zz_late1_IntAluPlugin_logic_alu_result_5 = execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
  assign _zz_late1_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_late1_IntAluPlugin_logic_alu_result_5};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[4 : 0];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[0],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[1],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[2],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[3],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[4],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[5],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[6],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[7],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[8],{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_2,_zz_late1_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_late1_BarrelShifterPlugin_logic_shift_shifted_1) >>> late1_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_late1_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1 && execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]),late1_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched = {late1_BarrelShifterPlugin_logic_shift_shifted[0],{late1_BarrelShifterPlugin_logic_shift_shifted[1],{late1_BarrelShifterPlugin_logic_shift_shifted[2],{late1_BarrelShifterPlugin_logic_shift_shifted[3],{late1_BarrelShifterPlugin_logic_shift_shifted[4],{late1_BarrelShifterPlugin_logic_shift_shifted[5],{late1_BarrelShifterPlugin_logic_shift_shifted[6],{late1_BarrelShifterPlugin_logic_shift_shifted[7],{late1_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_late1_BarrelShifterPlugin_logic_shift_patched_1,{_zz_late1_BarrelShifterPlugin_logic_shift_patched_2,_zz_late1_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_when_1 = (_zz_39 & (~ _zz_when_2));
  assign _zz_when_2 = (_zz_39 - 2'b01);
  assign _zz_FetchL1Plugin_logic_bus_cmd_payload_io = ((_zz_FetchL1Plugin_logic_bus_cmd_payload_address ? FetchL1Plugin_logic_refill_slots_0_isIo : 1'b0) | (_zz_FetchL1Plugin_logic_bus_cmd_payload_id ? FetchL1Plugin_logic_refill_slots_1_isIo : 1'b0));
  assign _zz_FetchL1Plugin_logic_ctrl_dataAccessFault = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error : 1'b0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error : 1'b0));
  assign _zz_FetchL1Plugin_logic_plru_write_payload_data_0 = 1'b0;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2 = fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2[1:0];
  assign _zz_BtbPlugin_logic_ras_ptr_push = (BtbPlugin_logic_ras_ptr_push + _zz_BtbPlugin_logic_ras_ptr_push_1);
  assign _zz_BtbPlugin_logic_ras_ptr_push_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_2};
  assign _zz_BtbPlugin_logic_ras_ptr_push_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_4};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue = (BtbPlugin_logic_ras_ptr_pop + _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1);
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4};
  assign _zz_WhiteboxerPlugin_logic_decodes_0_pc = {32'd0, decode_ctrls_0_down_PC_0};
  assign _zz_WhiteboxerPlugin_logic_decodes_1_pc = {32'd0, decode_ctrls_0_down_PC_1};
  assign _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = (|((FetchL1Plugin_pmaBuilder_addressBits & 32'h0) == 32'h0));
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault);
  assign _zz_FetchL1WishbonePlugin_logic_bus_ADR = (FetchL1Plugin_logic_bus_cmd_payload_address >>> 3'd6);
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_Decode_UOP_lane0[31 : 20];
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 25],execute_ctrl1_down_Decode_UOP_lane0[11 : 7]};
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) + $signed(early0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1 = _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3 = execute_ctrl2_down_SrcStageables_REVERT_lane0;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2 = {31'd0, _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz__zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = execute_ctrl3_down_Decode_UOP_lane0[31 : 20];
  assign _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 = ($signed(execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0) + $signed(late0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1 = _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3 = execute_ctrl4_down_SrcStageables_REVERT_lane0;
  assign _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2 = {31'd0, _zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz__zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = execute_ctrl1_down_Decode_UOP_lane1[31 : 20];
  assign _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 = ($signed(execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1) + $signed(early1_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1 = _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2;
  assign _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3 = execute_ctrl2_down_SrcStageables_REVERT_lane1;
  assign _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2 = {31'd0, _zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3};
  assign _zz__zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = execute_ctrl3_down_Decode_UOP_lane1[31 : 20];
  assign _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 = ($signed(execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1) + $signed(late1_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1 = _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2;
  assign _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3 = execute_ctrl4_down_SrcStageables_REVERT_lane1;
  assign _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2 = {31'd0, _zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3};
  assign _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent_1 = FpuAddPlugin_logic_addPort_cmd_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent = {{1{_zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent_1[11]}}, _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent_1};
  assign _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent = FpuMulPlugin_logic_addPort_cmd_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent = FpuAddPlugin_logic_addPort_cmd_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent = FpuMulPlugin_logic_addPort_cmd_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent_1[12 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent_1 = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1[16 : 4];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1[121 : 17];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent_1[11 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent_1 = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1[15 : 4];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1[67 : 16];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21 = _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_1 = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_2) - $signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_4));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_3 = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_2 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_3[11]}}, _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_3};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21_4 = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12 = _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_1 = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_2) - $signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_3));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_2 = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_4 = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_3 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_4[11]}}, _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12_4};
  assign _zz__zz_when_AFix_l1168 = FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12;
  assign _zz__zz_when_AFix_l1168_1 = FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_2 = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_1 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_2[11]}}, _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_2};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger = ({53'd0,FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa} <<< 6'd53);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa = (_zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_1 + _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_4);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_2 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger ? FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mantissa : _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_3);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_1 = {1'd0, _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_2};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_3 = ({53'd0,FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mantissa} <<< 6'd53);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa_4 = ({105'd0,1'b1} <<< 7'd105);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted = (_zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_1 + _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_4);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_2 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger ? _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_3 : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mantissa);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_1 = {1'd0, _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_2};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_3 = ({53'd0,FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mantissa} <<< 6'd53);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted_4 = ({105'd0,1'b1} <<< 7'd105);
  assign _zz__zz_when_Utils_l1585_13 = (_zz_when_Utils_l1585_14 >>> 1'b1);
  assign _zz__zz_when_Utils_l1585_12 = (_zz_when_Utils_l1585_13 >>> 2'b10);
  assign _zz__zz_when_Utils_l1585_11 = (_zz_when_Utils_l1585_12 >>> 3'b100);
  assign _zz__zz_when_Utils_l1585_10 = (_zz_when_Utils_l1585_11 >>> 4'b1000);
  assign _zz__zz_when_Utils_l1585_9 = (_zz_when_Utils_l1585_10 >>> 5'h10);
  assign _zz__zz_when_Utils_l1585_8 = (_zz_when_Utils_l1585_9 >>> 6'h20);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter = (_zz_when_Utils_l1585_8 >>> 7'h40);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_3 = _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_2 = {107'd0, _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_3};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger ? FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent : _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_1);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_2 = FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_1 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_2[11]}}, _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent_2};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_1 = _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_2;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_2 = _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_3;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_3 = ({FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_needSub,(FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_needSub ? (~ _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned) : _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned)} + _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_4);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_5 = (FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_needSub && (! FpuAddSharedPlugin_logic_pip_node_2_adder_math_roundingScrap));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_4 = {107'd0, _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_5};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa = _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_1 = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_2) + $signed(_zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_5));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_3 = {1'b0,_zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_4};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_2 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_3[107]}}, _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_3};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_4 = ({1'd0,FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xMantissa} <<< 1'd1);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_6 = FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_5 = {{1{_zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_6[107]}}, _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa_6};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_1 = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_2) + $signed(_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_7));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_2 = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_3;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_3 = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_4) - $signed(_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_5));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_4 = FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_6 = {1'b0,FpuAddSharedPlugin_logic_pip_node_4_adder_norm_shift};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_5 = {{5{_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_6[7]}}, _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_6};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_8 = {1'b0,1'b1};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_7 = {{11{_zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_8[1]}}, _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent_8};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa = {FpuAddSharedPlugin_logic_pip_node_4_adder_result_mantissa,FpuAddSharedPlugin_logic_pip_node_4_adder_math_roundingScrap};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent_1;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent_1 = FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent;
  assign _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_exponent = FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent = FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent = FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent = FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent = FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent = FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent = FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent = FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_exponent = FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_exponent = FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent = FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent;
  assign _zz_execute_ctrl2_down_MUL_SRC1_lane0_1 = {(execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_up_integer_RS1_lane0[31]),execute_ctrl2_up_integer_RS1_lane0};
  assign _zz_execute_ctrl2_down_MUL_SRC1_lane0 = {{21{_zz_execute_ctrl2_down_MUL_SRC1_lane0_1[32]}}, _zz_execute_ctrl2_down_MUL_SRC1_lane0_1};
  assign _zz_execute_ctrl2_down_MUL_SRC2_lane0_1 = {(execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_up_integer_RS2_lane0[31]),execute_ctrl2_up_integer_RS2_lane0};
  assign _zz_execute_ctrl2_down_MUL_SRC2_lane0 = {{21{_zz_execute_ctrl2_down_MUL_SRC2_lane0_1[32]}}, _zz_execute_ctrl2_down_MUL_SRC2_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = {{36{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = {{36{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = {{19{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[33 : 17]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = {{19{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = {{2{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[50 : 34]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = {{2{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1[20]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_1 = execute_ctrl2_down_MUL_SRC1_lane0[53 : 51];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0_2 = execute_ctrl2_down_MUL_SRC2_lane0[53 : 51];
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_8 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_9 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_10 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_11 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_12 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_13 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_15 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_16 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_17 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_18 = {3'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6};
  assign _zz_early0_DivPlugin_logic_processing_selected = early0_DivPlugin_logic_processing_div_io_rsp_payload_remain[31:0];
  assign _zz_early0_DivPlugin_logic_processing_selected_1 = early0_DivPlugin_logic_processing_div_io_rsp_payload_result[31:0];
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1 = ((early0_DivPlugin_logic_processing_divRevertResult ? (~ _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) : _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) + _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3 = early0_DivPlugin_logic_processing_divRevertResult;
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2 = {31'd0, _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3};
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_code = {2'd0, early0_EnvPlugin_logic_exe_privilege};
  assign _zz_early0_BranchPlugin_pcCalc_target_b = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[19 : 12]},execute_ctrl2_down_Decode_UOP_lane0[20]},execute_ctrl2_down_Decode_UOP_lane0[30 : 21]},1'b0};
  assign _zz_early0_BranchPlugin_pcCalc_target_b_1 = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign _zz_early0_BranchPlugin_pcCalc_target_b_2 = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[7]},execute_ctrl2_down_Decode_UOP_lane0[30 : 25]},execute_ctrl2_down_Decode_UOP_lane0[11 : 8]},1'b0};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = ($signed(early0_BranchPlugin_pcCalc_target_a) + $signed(early0_BranchPlugin_pcCalc_target_b));
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1 = ({1'd0,early0_BranchPlugin_pcCalc_slices} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = {29'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1 = ({1'd0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = {30'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1};
  assign _zz_early1_BranchPlugin_pcCalc_target_b = {{{{execute_ctrl2_down_Decode_UOP_lane1[31],execute_ctrl2_down_Decode_UOP_lane1[19 : 12]},execute_ctrl2_down_Decode_UOP_lane1[20]},execute_ctrl2_down_Decode_UOP_lane1[30 : 21]},1'b0};
  assign _zz_early1_BranchPlugin_pcCalc_target_b_1 = execute_ctrl2_down_Decode_UOP_lane1[31 : 20];
  assign _zz_early1_BranchPlugin_pcCalc_target_b_2 = {{{{execute_ctrl2_down_Decode_UOP_lane1[31],execute_ctrl2_down_Decode_UOP_lane1[7]},execute_ctrl2_down_Decode_UOP_lane1[30 : 25]},execute_ctrl2_down_Decode_UOP_lane1[11 : 8]},1'b0};
  assign _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = ($signed(early1_BranchPlugin_pcCalc_target_a) + $signed(early1_BranchPlugin_pcCalc_target_b));
  assign _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1 = ({1'd0,early1_BranchPlugin_pcCalc_slices} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = {29'd0, _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1};
  assign _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1 = ({1'd0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1} <<< 1'd1);
  assign _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = {30'd0, _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1};
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = (4'b0001 <<< fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign _zz_AlignerPlugin_logic_extractors_0_redo_8 = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? _zz_AlignerPlugin_logic_extractors_0_redo_9 : _zz_AlignerPlugin_logic_extractors_0_redo_10) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? _zz_AlignerPlugin_logic_extractors_0_redo_11 : _zz_AlignerPlugin_logic_extractors_0_redo_12)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? _zz_AlignerPlugin_logic_extractors_0_redo_13 : _zz_AlignerPlugin_logic_extractors_0_redo_14) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? _zz_AlignerPlugin_logic_extractors_0_redo_15 : _zz_AlignerPlugin_logic_extractors_0_redo_16))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? _zz_AlignerPlugin_logic_extractors_0_redo_17 : _zz_AlignerPlugin_logic_extractors_0_redo_18) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? _zz_AlignerPlugin_logic_extractors_0_redo_19 : _zz_AlignerPlugin_logic_extractors_0_redo_20)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? _zz_AlignerPlugin_logic_extractors_0_redo_21 : _zz_AlignerPlugin_logic_extractors_0_redo_22) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? _zz_AlignerPlugin_logic_extractors_0_redo_23 : _zz_AlignerPlugin_logic_extractors_0_redo_24))));
  assign _zz_AlignerPlugin_logic_extractors_1_redo_7 = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? _zz_AlignerPlugin_logic_extractors_1_redo_8 : _zz_AlignerPlugin_logic_extractors_1_redo_9) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? _zz_AlignerPlugin_logic_extractors_1_redo_10 : _zz_AlignerPlugin_logic_extractors_1_redo_11)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? _zz_AlignerPlugin_logic_extractors_1_redo_12 : _zz_AlignerPlugin_logic_extractors_1_redo_13) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? _zz_AlignerPlugin_logic_extractors_1_redo_14 : _zz_AlignerPlugin_logic_extractors_1_redo_15))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? _zz_AlignerPlugin_logic_extractors_1_redo_16 : _zz_AlignerPlugin_logic_extractors_1_redo_17) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? _zz_AlignerPlugin_logic_extractors_1_redo_18 : _zz_AlignerPlugin_logic_extractors_1_redo_19)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? AlignerPlugin_logic_scanners_7_redo : 1'b0)));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26 = {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},12'h0};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 = {6'd0, _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35 = {{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36 = {{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_37 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_38 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_39 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_40 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[1]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice = {1'd0, decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26 = {{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},12'h0};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1 = {AlignerPlugin_logic_extractors_1_ctx_instruction[12],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 = {6'd0, _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35 = {{{3'b000,AlignerPlugin_logic_extractors_1_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36 = {{{3'b000,AlignerPlugin_logic_extractors_1_ctx_instruction[9 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_37 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_38 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_39 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_40 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4[1]};
  assign _zz_decode_ctrls_0_up_Decode_DOP_ID_1_1 = decode_ctrls_0_up_LANE_SEL_0;
  assign _zz_decode_ctrls_0_up_Decode_DOP_ID_1 = {9'd0, _zz_decode_ctrls_0_up_Decode_DOP_ID_1_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice = {1'd0, decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1};
  assign _zz_LsuPlugin_logic_storeBuffer_ops_popPtr_1 = LsuPlugin_logic_storeBuffer_ops_pip_node_0_isFiring;
  assign _zz_LsuPlugin_logic_storeBuffer_ops_popPtr = {5'd0, _zz_LsuPlugin_logic_storeBuffer_ops_popPtr_1};
  assign _zz__zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1 = _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address[4:0];
  assign _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr_1 = LsuPlugin_logic_storeBuffer_push_valid;
  assign _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr = {5'd0, _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr_1};
  assign _zz_LsuPlugin_logic_storeBuffer_ops_mem_port_1 = LsuPlugin_logic_storeBuffer_ops_pushPtr[4:0];
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId_1 = LsuPlugin_logic_onAddress0_ls_port_fire;
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId = {11'd0, _zz_LsuPlugin_logic_onAddress0_ls_storeId_1};
  assign _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address = ({6'd0,LsuPlugin_logic_flusher_cmdCounter} <<< 3'd6);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1 = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2 = execute_ctrl4_down_integer_RS2_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? (~ LsuPlugin_logic_onCtrl_rva_srcBuffer) : LsuPlugin_logic_onCtrl_rva_srcBuffer);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? 2'b01 : 2'b00);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4 = {{30{_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5[1]}}, _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5};
  assign _zz_LsuPlugin_logic_trapPort_payload_code = (execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 ? (execute_ctrl4_down_LsuL1_STORE_lane0 ? 3'b110 : 3'b100) : 3'b000);
  assign _zz_LsuPlugin_logic_flusher_cmdCounter = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign _zz_FpuPackerPlugin_logic_s0_remapped_1_exponent = FpuMulPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent_1 = FpuSqrtPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent = {{2{_zz_FpuPackerPlugin_logic_s0_remapped_2_exponent_1[10]}}, _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent_1};
  assign _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent_1 = FpuXxPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent = {{1{_zz_FpuPackerPlugin_logic_s0_remapped_3_exponent_1[11]}}, _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent_1};
  assign _zz_FpuPackerPlugin_logic_s0_remapped_4_exponent = FpuDivPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_FpuPackerPlugin_logic_s0_remapped_5_exponent = FpuAddSharedPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent_1[12 : 0];
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent_1 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1[16 : 4];
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1[70 : 17];
  assign _zz_65 = (_zz_66 + _zz_68);
  assign _zz_70 = {FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[4],FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[3]};
  assign _zz_69 = {1'd0, _zz_70};
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL = _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL_1;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL_1 = ((FpuPackerPlugin_logic_pip_node_0_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? 11'h401 : 11'h781);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE = FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_2 = FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_1 = {{2{_zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_2[10]}}, _zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_2};
  assign _zz__zz_when_AFix_l1168_1_1 = ($signed(_zz__zz_when_AFix_l1168_1_2) - $signed(_zz__zz_when_AFix_l1168_1_4));
  assign _zz__zz_when_AFix_l1168_1_3 = FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL;
  assign _zz__zz_when_AFix_l1168_1_2 = {{2{_zz__zz_when_AFix_l1168_1_3[10]}}, _zz__zz_when_AFix_l1168_1_3};
  assign _zz__zz_when_AFix_l1168_1_4 = FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  assign _zz__zz_when_Utils_l1585_7 = (_zz_when_Utils_l1585_15 >>> 1'b1);
  assign _zz__zz_when_Utils_l1585_6 = (_zz_when_Utils_l1585_7 >>> 2'b10);
  assign _zz__zz_when_Utils_l1585_5 = (_zz_when_Utils_l1585_6 >>> 3'b100);
  assign _zz__zz_when_Utils_l1585_4 = (_zz_when_Utils_l1585_5 >>> 4'b1000);
  assign _zz__zz_when_Utils_l1585_3 = (_zz_when_Utils_l1585_4 >>> 5'h10);
  assign _zz__zz_FpuPackerPlugin_logic_s1_subnormal_manShifter = (_zz_when_Utils_l1585_3 >>> 6'h20);
  assign _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_2 = (_zz_FpuPackerPlugin_logic_s1_subnormal_manShifter | _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_3);
  assign _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_4 = _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1;
  assign _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_3 = {54'd0, _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_4};
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted_1 = (|FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED[28 : 0]);
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted = {1'd0, _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted_1};
  assign _zz_FpuPackerPlugin_logic_s1_incrBy = ({29'd0,1'b1} <<< 5'd29);
  assign _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry = (FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED >>> 2'd2);
  assign _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_2 = {1'b0,FpuPackerPlugin_logic_s1_incrBy};
  assign _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_1 = {22'd0, _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_2};
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR = _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_1;
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_1 = ($signed(_zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_2) + $signed(_zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_3));
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_2 = FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_4 = {1'b0,FpuPackerPlugin_logic_s1_MAN_CARRY};
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_3 = {{11{_zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_4[1]}}, _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR_4};
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT = (FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR ? FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR : _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT_1);
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT_1 = FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT = (FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED >>> 2'd2);
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL = _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_1;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_1 = ($signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_2) - $signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_4));
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_3 = FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_2 = {{2{_zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_3[10]}}, _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_3};
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL_4 = FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP = ((! FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL) ? _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_1 : 13'h0);
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_1 = ($signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_2) - $signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_3));
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_2 = FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_4 = FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_3 = {{2{_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_4[10]}}, _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_4};
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX = _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX_1;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX_1 = ((FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? 11'h3ff : 11'h07f);
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN = _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN_1;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN_1 = ((FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? 12'hbcc : 12'hf69);
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_1 = FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW = {{2{_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_1[10]}}, _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_1};
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_2 = FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW = FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_2 = FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_1 = {{1{_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_2[11]}}, _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_2};
  assign _zz_FpuPackerPlugin_logic_s2_fwb_value = FpuPackerPlugin_logic_pip_node_2_s2_EXP[10:0];
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent = FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL = FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s0_VALUE_exponent = FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL = FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL;
  assign _zz_FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT = FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT;
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = {early0_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[0]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = {early0_BranchPlugin_logic_jumpLogic_history_shifter_1,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[1]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_3 = {early0_BranchPlugin_logic_jumpLogic_history_shifter_2,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[2]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_4 = {early0_BranchPlugin_logic_jumpLogic_history_shifter_3,execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_1 = {early1_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[0]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_2 = {early1_BranchPlugin_logic_jumpLogic_history_shifter_1,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[1]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_3 = {early1_BranchPlugin_logic_jumpLogic_history_shifter_2,execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[2]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_4 = {early1_BranchPlugin_logic_jumpLogic_history_shifter_3,execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1};
  assign _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED = _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_1;
  assign _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_1 = (PrefetcherRptPlugin_logic_pip_node_1_PROBE_address - _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_2);
  assign _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED_2 = {16'd0, PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address};
  assign _zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK = ((_zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK_1 ^ PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address) >>> 3'd6);
  assign _zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK_1 = PrefetcherRptPlugin_logic_pip_node_1_PROBE_address[15:0];
  assign _zz__zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT = PrefetcherRptPlugin_logic_pip_node_2_STRIDE_EXTENDED[15 : 12];
  assign _zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT_1 = PrefetcherRptPlugin_logic_pip_node_2_STRIDE_EXTENDED[11:0];
  assign _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed_1 = {1'b0,PrefetcherRptPlugin_logic_pip_node_2_NEW_BLOCK};
  assign _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed = {2'd0, _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed_1};
  assign _zz__zz_when_UInt_l128_1_1 = {1'b0,2'b11};
  assign _zz__zz_when_UInt_l128_1 = {3'd0, _zz__zz_when_UInt_l128_1_1};
  assign _zz_PrefetcherRptPlugin_logic_storage_write_payload_data_address = PrefetcherRptPlugin_logic_pip_node_2_PROBE_address[15:0];
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_1 = ((PrefetcherRptPlugin_logic_onCtrl_advanceAllowed < _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_2) ? PrefetcherRptPlugin_logic_onCtrl_advanceAllowed : _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_3);
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_2 = {2'd0, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to};
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_3 = {2'd0, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to};
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_2 = (($signed(PrefetcherRptPlugin_logic_pip_node_2_STRIDE) < $signed(_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_3)) ? PrefetcherRptPlugin_logic_pip_node_2_STRIDE : _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_4);
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_3 = {{5{_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride[6]}}, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride};
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_4 = {{5{_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride[6]}}, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride};
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_5 = (($signed(PrefetcherRptPlugin_logic_pip_node_2_STRIDE) < $signed(_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_6)) ? _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_7 : PrefetcherRptPlugin_logic_pip_node_2_STRIDE);
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_6 = {{4{_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1[7]}}, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1};
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_7 = {{4{_zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1[7]}}, _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1};
  assign _zz_when_Prefetcher_l216 = {2'd0, PrefetcherRptPlugin_logic_onCtrl_advanceSubed};
  assign _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io_1 = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = (|((LsuPlugin_pmaBuilder_io_addressBits & 32'h0) == 32'h0));
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io = (|_zz_LsuPlugin_logic_onPma_io_rsp_fault);
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_1 = {late0_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[0]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_2 = {late0_BranchPlugin_logic_jumpLogic_history_shifter_1,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[1]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_3 = {late0_BranchPlugin_logic_jumpLogic_history_shifter_2,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[2]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_4 = {late0_BranchPlugin_logic_jumpLogic_history_shifter_3,execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_1 = {late1_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[0]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_2 = {late1_BranchPlugin_logic_jumpLogic_history_shifter_1,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[1]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_3 = {late1_BranchPlugin_logic_jumpLogic_history_shifter_2,execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[2]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_4 = {late1_BranchPlugin_logic_jumpLogic_history_shifter_3,execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1};
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0 = (|{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000044) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000018) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS1_ENABLE_0_1) == 32'h00002000),{(_zz_decode_ctrls_1_down_RS1_ENABLE_0_2 == _zz_decode_ctrls_1_down_RS1_ENABLE_0_3),(_zz_decode_ctrls_1_down_RS1_ENABLE_0_4 == _zz_decode_ctrls_1_down_RS1_ENABLE_0_5)}}}}});
  assign _zz_decode_ctrls_1_down_RS1_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[19 : 15];
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000034) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h40000060) == 32'h00000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS2_ENABLE_0_1) == 32'h00000020),{(_zz_decode_ctrls_1_down_RS2_ENABLE_0_2 == _zz_decode_ctrls_1_down_RS2_ENABLE_0_3),{_zz_decode_ctrls_1_down_RS2_ENABLE_0_4,_zz_decode_ctrls_1_down_RS2_ENABLE_0_5}}}}}});
  assign _zz_decode_ctrls_1_down_RS2_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[24 : 20];
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000048) == 32'h00000048),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001010) == 32'h00001010),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002008) == 32'h00002008),{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0,{(_zz_decode_ctrls_1_down_RD_ENABLE_0_1 == _zz_decode_ctrls_1_down_RD_ENABLE_0_2),{_zz_decode_ctrls_1_down_RD_ENABLE_0_3,{_zz_decode_ctrls_1_down_RD_ENABLE_0_4,_zz_decode_ctrls_1_down_RD_ENABLE_0_5}}}}}}}});
  assign _zz_decode_ctrls_1_down_RD_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7];
  assign _zz_decode_ctrls_1_down_RS3_ENABLE_0 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0);
  assign _zz_decode_ctrls_1_down_RS3_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[31 : 27];
  assign _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1 = ((! decode_ctrls_1_down_Prediction_ALIGN_REDO_0) ? _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = {30'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1};
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 = ({1'd0,decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0} <<< 1'd1);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1 = (|{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000044) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000018) == 32'h0),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_RS1_ENABLE_1_1) == 32'h00002000),{(_zz_decode_ctrls_1_down_RS1_ENABLE_1_2 == _zz_decode_ctrls_1_down_RS1_ENABLE_1_3),(_zz_decode_ctrls_1_down_RS1_ENABLE_1_4 == _zz_decode_ctrls_1_down_RS1_ENABLE_1_5)}}}}});
  assign _zz_decode_ctrls_1_down_RS1_PHYS_1 = decode_ctrls_1_down_Decode_INSTRUCTION_1[19 : 15];
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000034) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h40000060) == 32'h00000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_RS2_ENABLE_1_1) == 32'h00000020),{(_zz_decode_ctrls_1_down_RS2_ENABLE_1_2 == _zz_decode_ctrls_1_down_RS2_ENABLE_1_3),{_zz_decode_ctrls_1_down_RS2_ENABLE_1_4,_zz_decode_ctrls_1_down_RS2_ENABLE_1_5}}}}}});
  assign _zz_decode_ctrls_1_down_RS2_PHYS_1 = decode_ctrls_1_down_Decode_INSTRUCTION_1[24 : 20];
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000048) == 32'h00000048),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001010) == 32'h00001010),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002008) == 32'h00002008),{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1,{(_zz_decode_ctrls_1_down_RD_ENABLE_1_1 == _zz_decode_ctrls_1_down_RD_ENABLE_1_2),{_zz_decode_ctrls_1_down_RD_ENABLE_1_3,{_zz_decode_ctrls_1_down_RD_ENABLE_1_4,_zz_decode_ctrls_1_down_RD_ENABLE_1_5}}}}}}}});
  assign _zz_decode_ctrls_1_down_RD_PHYS_1 = decode_ctrls_1_down_Decode_INSTRUCTION_1[11 : 7];
  assign _zz_decode_ctrls_1_down_RS3_ENABLE_1 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1);
  assign _zz_decode_ctrls_1_down_RS3_PHYS_1 = decode_ctrls_1_down_Decode_INSTRUCTION_1[31 : 27];
  assign _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4 = ((! decode_ctrls_1_down_Prediction_ALIGN_REDO_1) ? _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3 = {30'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4};
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5 = ({1'd0,decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1} <<< 1'd1);
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = LearnPlugin_logic_learn_payload_history;
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash_2[1:0];
  assign _zz_BtbPlugin_logic_memWrite_payload_address = (LearnPlugin_logic_learn_payload_pcOnLastSlice >>> 2'd3);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent = (FpuUnpack_RS1_f64_exponent - 11'h3ff);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa = ({29'd0,FpuUnpack_RS1_f32_mantissa} <<< 5'd29);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_1 = (_zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_2 - 11'h07f);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_2 = {3'd0, FpuUnpack_RS1_f32_exponent};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_1 = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent = {{1{_zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_1[10]}}, _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_1};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_2 = FpuUnpack_RS1_normalizer_exponent;
  assign _zz_FpuUnpack_RS1_normalizer_exponent = ($signed(FpuUnpack_RS1_recodedExpSub) - $signed(_zz_FpuUnpack_RS1_normalizer_exponent_1));
  assign _zz_FpuUnpack_RS1_normalizer_exponent_2 = {1'b0,FpuUnpackerPlugin_logic_unpacker_results_0_payload_shift};
  assign _zz_FpuUnpack_RS1_normalizer_exponent_1 = {{5{_zz_FpuUnpack_RS1_normalizer_exponent_2[6]}}, _zz_FpuUnpack_RS1_normalizer_exponent_2};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent = (FpuUnpack_RS2_f64_exponent - 11'h3ff);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa = ({29'd0,FpuUnpack_RS2_f32_mantissa} <<< 5'd29);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_1 = (_zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_2 - 11'h07f);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_2 = {3'd0, FpuUnpack_RS2_f32_exponent};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_1 = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent = {{1{_zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_1[10]}}, _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_1};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_2 = FpuUnpack_RS2_normalizer_exponent;
  assign _zz_FpuUnpack_RS2_normalizer_exponent = ($signed(FpuUnpack_RS2_recodedExpSub) - $signed(_zz_FpuUnpack_RS2_normalizer_exponent_1));
  assign _zz_FpuUnpack_RS2_normalizer_exponent_2 = {1'b0,FpuUnpackerPlugin_logic_unpacker_results_0_payload_shift};
  assign _zz_FpuUnpack_RS2_normalizer_exponent_1 = {{5{_zz_FpuUnpack_RS2_normalizer_exponent_2[6]}}, _zz_FpuUnpack_RS2_normalizer_exponent_2};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent = (FpuUnpack_RS3_f64_exponent - 11'h3ff);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa = ({29'd0,FpuUnpack_RS3_f32_mantissa} <<< 5'd29);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_1 = (_zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_2 - 11'h07f);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_2 = {3'd0, FpuUnpack_RS3_f32_exponent};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_1 = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent = {{1{_zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_1[10]}}, _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_1};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_2 = FpuUnpack_RS3_normalizer_exponent;
  assign _zz_FpuUnpack_RS3_normalizer_exponent = ($signed(FpuUnpack_RS3_recodedExpSub) - $signed(_zz_FpuUnpack_RS3_normalizer_exponent_1));
  assign _zz_FpuUnpack_RS3_normalizer_exponent_2 = {1'b0,FpuUnpackerPlugin_logic_unpacker_results_0_payload_shift};
  assign _zz_FpuUnpack_RS3_normalizer_exponent_1 = {{5{_zz_FpuUnpack_RS3_normalizer_exponent_2[6]}}, _zz_FpuUnpack_RS3_normalizer_exponent_2};
  assign _zz_io_inputs_1_payload_data = execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  assign _zz_FpuUnpackerPlugin_logic_packPort_cmd_value_exponent = (6'h34 - FpuUnpackerPlugin_logic_onCvt_fsmResult_shift);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_2[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_2 = (|{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005c) == 32'h00000004),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffe02050) == 32'h00202050),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffe01050) == 32'h00201050),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_3) == 32'h00102050),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_4) == 32'h00101050)}}}}});
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h90000060) == 32'h10000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h60000060) == 32'h00000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h22000060) == 32'h00000040),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hb0000060) == 32'h80000040)}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_4}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_15,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_14,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_3}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_16 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_17[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_17 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_15,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_14,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_18,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_19}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000060) == 32'h00000060),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000030) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001050) == 32'h00001000),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000058) == 32'h0)}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h18000050) == 32'h18000050),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hb0000050) == 32'h90000050)}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0_1[0];
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0_1 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_2[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_2 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0_1 = (|((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h98000070) == 32'h10000050));
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0_1[0];
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0_1 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_2[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_2 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h18000070) == 32'h18000050),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hb0000070) == 32'h90000050)});
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0_1 = (|((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hd0000070) == 32'h40000050));
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_2[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_2 = (|{_zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000005c) == 32'h00000004),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffe02050) == 32'h00202050),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffe01050) == 32'h00201050),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_3) == 32'h00102050),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_4) == 32'h00101050)}}}}});
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h90000060) == 32'h10000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h60000060) == 32'h00000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h22000060) == 32'h00000040),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hb0000060) == 32'h80000040)}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_4}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_15,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_14,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_3}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_16 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_17[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_17 = (|{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_15,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_13,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_14,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_12,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_11,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_10,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_9,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_8,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_7,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_18,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_19}}}}}}}}}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000060) == 32'h00000060),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000030) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001050) == 32'h00001000),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000058) == 32'h0)}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1,{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h18000050) == 32'h18000050),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hb0000050) == 32'h90000050)}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1_1[0];
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1_1 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_2[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_2 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1_1 = (|((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h98000070) == 32'h10000050));
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1_1[0];
  assign _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1_1 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_2[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_2 = (|_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h18000070) == 32'h18000050),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hb0000070) == 32'h90000050)});
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1_1 = (|((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hd0000070) == 32'h40000050));
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0 = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0_1 = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0 = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0_1 = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_FpuCmpPlugin_logic_iwb_payload = execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0 = _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_1;
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_1 = ($signed(_zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_2) - $signed(_zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_4));
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_3 = {1'b0,5'h1f};
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_2 = {{6{_zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_3[5]}}, _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_3};
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0_4 = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz__zz_when_Utils_l1585_2 = (_zz_when_Utils_l1585_16 >>> 1'b1);
  assign _zz__zz_when_Utils_l1585_1 = (_zz_when_Utils_l1585_2 >>> 2'b10);
  assign _zz__zz_when_Utils_l1585 = (_zz_when_Utils_l1585_1 >>> 3'b100);
  assign _zz__zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 = (_zz_when_Utils_l1585 >>> 4'b1000);
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 = _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1;
  assign _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 = {53'd0, _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3};
  assign _zz__zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 >>> 3'd4);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 >>> 1'b1);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 >>> 2'b10);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 >>> 3'b100);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 >>> 4'b1000);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4 >>> 5'h10);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6_1 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5 >>> 6'h20);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_2 = _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_1 = {53'd0, _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_2};
  assign _zz_FpuF2iPlugin_logic_onResult_inverter = {31'd0, execute_ctrl4_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0};
  assign _zz_FpuF2iPlugin_logic_onResult_expMax_1 = ((FpuF2iPlugin_logic_onResult_i64 ? 6'h3e : _zz_FpuF2iPlugin_logic_onResult_expMax_2) + _zz_FpuF2iPlugin_logic_onResult_expMax_4);
  assign _zz_FpuF2iPlugin_logic_onResult_expMax_3 = 5'h1e;
  assign _zz_FpuF2iPlugin_logic_onResult_expMax_2 = {1'd0, _zz_FpuF2iPlugin_logic_onResult_expMax_3};
  assign _zz_FpuF2iPlugin_logic_onResult_expMax_5 = _zz_FpuF2iPlugin_logic_onResult_expMax;
  assign _zz_FpuF2iPlugin_logic_onResult_expMax_4 = {5'd0, _zz_FpuF2iPlugin_logic_onResult_expMax_5};
  assign _zz_FpuF2iPlugin_logic_onResult_expMin_1 = 5'h1f;
  assign _zz_FpuF2iPlugin_logic_onResult_expMin = {1'd0, _zz_FpuF2iPlugin_logic_onResult_expMin_1};
  assign _zz_FpuF2iPlugin_logic_onResult_overflow_1 = {1'b0,FpuF2iPlugin_logic_onResult_expMax};
  assign _zz_FpuF2iPlugin_logic_onResult_overflow = {{5{_zz_FpuF2iPlugin_logic_onResult_overflow_1[6]}}, _zz_FpuF2iPlugin_logic_onResult_overflow_1};
  assign _zz_FpuF2iPlugin_logic_onResult_overflow_2 = execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_FpuF2iPlugin_logic_onResult_underflow_1 = {1'b0,FpuF2iPlugin_logic_onResult_expMin};
  assign _zz_FpuF2iPlugin_logic_onResult_underflow = {{5{_zz_FpuF2iPlugin_logic_onResult_underflow_1[6]}}, _zz_FpuF2iPlugin_logic_onResult_underflow_1};
  assign _zz_FpuF2iPlugin_logic_onResult_underflow_2 = execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_FpuF2iPlugin_logic_onResult_underflow_3 = execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_FpuF2iPlugin_logic_onResult_underflow_5 = {1'b0,FpuF2iPlugin_logic_onResult_expMin};
  assign _zz_FpuF2iPlugin_logic_onResult_underflow_4 = {{5{_zz_FpuF2iPlugin_logic_onResult_underflow_5[6]}}, _zz_FpuF2iPlugin_logic_onResult_underflow_5};
  assign _zz_FpuAddPlugin_logic_addPort_cmd_rs1_exponent = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_FpuAddPlugin_logic_addPort_cmd_rs2_exponent = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_1;
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_1 = ($signed(_zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_2) + $signed(_zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_4));
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_3 = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_2 = {{1{_zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_3[11]}}, _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_3};
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_5 = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_4 = {{1{_zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_5[11]}}, _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0_5};
  assign _zz_execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0 = execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0 = _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_1;
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_1 = ($signed(_zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_2) + $signed(_zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_3));
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_2 = execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_4 = {1'b0,FpuMulPlugin_logic_norm_needShift};
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_3 = {{11{_zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_4[1]}}, _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0_4};
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0 = ({1'd0,execute_ctrl5_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0[103 : 0]} <<< 1'd1);
  assign _zz_FpuMulPlugin_logic_packPort_cmd_value_exponent = execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0;
  assign _zz_FpuMulPlugin_logic_addPort_cmd_rs1_exponent = execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0;
  assign _zz_FpuMulPlugin_logic_addPort_cmd_rs2_exponent = execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_FpuSqrtPlugin_logic_packPort_cmd_value_exponent = FpuSqrtPlugin_logic_onExecute_exp;
  assign _zz_FpuXxPlugin_logic_packPort_cmd_value_exponent = execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_early0_DivPlugin_logic_processing_a = {1'b1,execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa};
  assign _zz_early0_DivPlugin_logic_processing_b = {1'b1,execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa};
  assign _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0_1 = ((|early0_DivPlugin_logic_processing_div_io_rsp_payload_remain) || (|early0_DivPlugin_logic_processing_div_io_rsp_payload_result[0 : 0]));
  assign _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0 = {55'd0, _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0_1};
  assign _zz_FpuDivPlugin_logic_onExecute_mantissa_1 = execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0[0];
  assign _zz_FpuDivPlugin_logic_onExecute_mantissa = {53'd0, _zz_FpuDivPlugin_logic_onExecute_mantissa_1};
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent = _zz__zz_FpuDivPlugin_logic_onExecute_exponent_1;
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent_1 = ($signed(_zz__zz_FpuDivPlugin_logic_onExecute_exponent_2) - $signed(_zz__zz_FpuDivPlugin_logic_onExecute_exponent_4));
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent_3 = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent_2 = {{1{_zz__zz_FpuDivPlugin_logic_onExecute_exponent_3[11]}}, _zz__zz_FpuDivPlugin_logic_onExecute_exponent_3};
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent_5 = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz__zz_FpuDivPlugin_logic_onExecute_exponent_4 = {{1{_zz__zz_FpuDivPlugin_logic_onExecute_exponent_5[11]}}, _zz__zz_FpuDivPlugin_logic_onExecute_exponent_5};
  assign _zz_FpuDivPlugin_logic_onExecute_exponent_1 = ($signed(_zz_FpuDivPlugin_logic_onExecute_exponent_2) - $signed(_zz_FpuDivPlugin_logic_onExecute_exponent_3));
  assign _zz_FpuDivPlugin_logic_onExecute_exponent_2 = _zz_FpuDivPlugin_logic_onExecute_exponent;
  assign _zz_FpuDivPlugin_logic_onExecute_exponent_4 = {1'b0,FpuDivPlugin_logic_onExecute_needShift};
  assign _zz_FpuDivPlugin_logic_onExecute_exponent_3 = {{11{_zz_FpuDivPlugin_logic_onExecute_exponent_4[1]}}, _zz_FpuDivPlugin_logic_onExecute_exponent_4};
  assign _zz_FpuDivPlugin_logic_packPort_cmd_value_exponent = FpuDivPlugin_logic_onExecute_exponent;
  assign _zz_BtbPlugin_logic_memWrite_payload_address_1 = (DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice >>> 2'd3);
  assign _zz_BtbPlugin_logic_memRead_cmd_payload = (fetch_logic_ctrls_0_down_Fetch_WORD_PC >>> 2'd3);
  assign _zz_BtbPlugin_logic_ras_write_payload_data = (BtbPlugin_logic_applyIt_rasLogic_pushPc + 32'h00000002);
  assign _zz_DispatchPlugin_logic_inserter_0_trap = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_execute_ctrl0_up_LANE_SEL_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_cancel : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_cancel : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_cancel : 1'b0));
  assign _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0));
  assign _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0));
  assign _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0));
  assign _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0));
  assign _zz_execute_ctrl0_up_TRAP_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_execute_ctrl0_up_RS1_ENABLE_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RS2_ENABLE_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RD_ENABLE_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RS3_ENABLE_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_DispatchPlugin_logic_inserter_1_trap = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_execute_ctrl0_up_LANE_SEL_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_cancel : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_cancel : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_cancel : 1'b0));
  assign _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0));
  assign _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 : 1'b0));
  assign _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 : 1'b0));
  assign _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0));
  assign _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0));
  assign _zz_execute_ctrl0_up_TRAP_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_execute_ctrl0_up_RS1_ENABLE_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RS2_ENABLE_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RD_ENABLE_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_RS3_ENABLE_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 : 1'b0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 : 1'b0));
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_slices = {1'd0, _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1};
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1 = ({1'd0,TrapPlugin_logic_harts_0_trap_fsm_jumpOffset} <<< 1'd1);
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget = {29'd0, _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1};
  assign _zz_PcPlugin_logic_harts_0_self_pc_1 = (PcPlugin_logic_harts_0_self_increment ? 4'b1000 : 4'b0000);
  assign _zz_PcPlugin_logic_harts_0_self_pc = {28'd0, _zz_PcPlugin_logic_harts_0_self_pc_1};
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault = ((((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? late0_BranchPlugin_logic_pcPort_payload_fault : 1'b0)) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? late1_BranchPlugin_logic_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_3 ? early0_BranchPlugin_logic_pcPort_payload_fault : 1'b0))) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_4 ? early1_BranchPlugin_logic_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_5 ? PcPlugin_logic_harts_0_self_flow_payload_fault : 1'b0)));
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_fault : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = ({1'd0,(REG_CSR_2047 ? PrefetcherRptPlugin_logic_csr_disable : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_3858) ? 6'h2e : 6'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mpie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mpp : 2'b00)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = {19'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = ({17'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mprv : 1'b0)} <<< 5'd17);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = {14'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = {17'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? PrivilegedPlugin_logic_harts_0_m_cause_interrupt : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? PrivilegedPlugin_logic_harts_0_m_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_meip : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_mtip : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_msip : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_meie : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_mtie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_msie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? FpuCsrPlugin_api_rm : 3'b000)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? {FpuCsrPlugin_api_flags_NV,{FpuCsrPlugin_api_flags_DZ,{FpuCsrPlugin_api_flags_OF,{FpuCsrPlugin_api_flags_UF,FpuCsrPlugin_api_flags_NX}}}} : 5'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 = {27'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 = (REG_CSR_2 ? FpuCsrPlugin_api_rm : 3'b000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 = {29'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47 = (REG_CSR_1 ? {FpuCsrPlugin_api_flags_NV,{FpuCsrPlugin_api_flags_DZ,{FpuCsrPlugin_api_flags_OF,{FpuCsrPlugin_api_flags_UF,FpuCsrPlugin_api_flags_NX}}}} : 5'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46 = {27'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47};
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = CsrAccessPlugin_logic_fsm_interface_uop[19 : 15];
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {27'd0, _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 3'b001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 2'b01);
  assign _zz_CsrRamPlugin_logic_flush_counter_1 = (! CsrRamPlugin_logic_flush_done);
  assign _zz_CsrRamPlugin_logic_flush_counter = {2'd0, _zz_CsrRamPlugin_logic_flush_counter_1};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_9,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_8,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_7,{((execute_lane0_logic_decoding_decodingBits & 33'h102002070) == 33'h100002030),{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_6,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_5,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_4,{_zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2,_zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_3}}}}}}}}});
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h100003074) == 33'h100001010),((execute_lane0_logic_decoding_decodingBits & 33'h102003054) == 33'h100001010)});
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10);
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h002004074) == 33'h002000030));
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_11,((execute_lane0_logic_decoding_decodingBits & 33'h000003070) == 33'h000000070)});
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h100000044) == 33'h000000004),{((execute_lane0_logic_decoding_decodingBits & 33'h100002040) == 33'h000002000),((execute_lane0_logic_decoding_decodingBits & 33'h100001040) == 33'h0)}});
  assign _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h100003044) == 33'h000001000));
  assign _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1 = _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2[0];
  assign _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2 = (|_zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_1});
  assign _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0 = _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0,{_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_1,_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0}}});
  assign _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h060003034) == 33'h060001010));
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0a0000070) == 33'h020000050));
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0c0000070) == 33'h080000050));
  assign _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0b0000070) == 33'h080000050));
  assign _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0 = _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h030203050) == 33'h030000050));
  assign _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0 = _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h070003050) == 33'h060000050));
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000003048) == 33'h000000008));
  assign _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h098000060) == 33'h010000040)});
  assign _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0d0000070) == 33'h050000050));
  assign _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h058000070) == 33'h018000050));
  assign _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0 = _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0b0000070) == 33'h090000050));
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2 = (|{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000000028) == 33'h000000028),{((execute_lane0_logic_decoding_decodingBits & 33'h000001030) == 33'h000001030),{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3) == 33'h000002030),{(_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4 == _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5),{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6,{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_7,_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_8}}}}}}});
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_3 = _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_4[0];
  assign _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_4 = (|{_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0,{_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_1,_zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0}}}}}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_3,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_11,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_15,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_14,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_13,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_12,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_9,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_8,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_7,{_zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_2,_zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_3}}}}}}}}}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_9[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_9 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0}}}}}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_4 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_5[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_5 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_3,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_1 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_2 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_1 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_2 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_16 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_17[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_17 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_11,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_15,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_14,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_13,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_12,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_9,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_8,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_7,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_18,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_19}}}}}}}}}}});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = (|{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1 = (|_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0);
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000000040) == 33'h000000040),{((execute_lane0_logic_decoding_decodingBits & 33'h040000034) == 33'h040000030),((execute_lane0_logic_decoding_decodingBits & 33'h000006014) == 33'h000002010)}});
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1 = (|{_zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h000000034) == 33'h000000034)});
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000004010) == 33'h0),((execute_lane0_logic_decoding_decodingBits & 33'h020000060) == 33'h000000040)});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,((execute_lane0_logic_decoding_decodingBits & 33'h102000068) == 33'h100000020)}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h100004020) == 33'h100004020),{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h100000060) == 33'h100000060),{((execute_lane0_logic_decoding_decodingBits & 33'h102000028) == 33'h100000020),{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,((execute_lane0_logic_decoding_decodingBits & 33'h1b0000010) == 33'h1a0000010)}}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1,{((execute_lane0_logic_decoding_decodingBits & 33'h080000010) == 33'h080000010),{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0,_zz_execute_ctrl1_down_BYPASSED_AT_6_lane0}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1,{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_1,_zz_execute_ctrl1_down_BYPASSED_AT_6_lane0}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_1 = _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_2[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_2 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1,{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_1,_zz_execute_ctrl1_down_BYPASSED_AT_6_lane0}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_2 = _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_3[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_3 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1,{_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h010000010) == 33'h010000010),_zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_1}}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_3 = _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_4[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_4 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2,_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1 = (|{_zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0,{_zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_2[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_2 = (|{_zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0,{_zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}});
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000002010) == 33'h000002000),((execute_lane0_logic_decoding_decodingBits & 33'h000005000) == 33'h000001000)});
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2 = (|_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h040000000) == 33'h040000000));
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1[0];
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1 = (|{_zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0,_zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0});
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1 = (|{_zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000100020) == 33'h0),((execute_lane0_logic_decoding_decodingBits & 33'h080006000) == 33'h0)}});
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000005000) == 33'h000004000),_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1[0];
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1 = (|_zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000004000) == 33'h000004000));
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1 = (|_zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1 = (|_zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0);
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_1 = _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_2[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_2 = (|_zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0);
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_1 = _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_2[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_2 = (|_zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0);
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_1 = _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_2[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h008002000) == 33'h0),_zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0});
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000001000) == 33'h0));
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000000028) == 33'h0),{((execute_lane0_logic_decoding_decodingBits & 33'h008002008) == 33'h000002008),((execute_lane0_logic_decoding_decodingBits & 33'h010002008) == 33'h000002008)}});
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h008000020) == 33'h008000020),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000000028) == 33'h000000020),((execute_lane0_logic_decoding_decodingBits & 33'h000206000) == 33'h000206000)}}});
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000002008) == 33'h000002008));
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_2 = (|_zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0);
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000006000) == 33'h000006000));
  assign _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0 = _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h008000000) == 33'h008000000));
  assign _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000000010) == 33'h0));
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_1 = _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_2[0];
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_2 = (|_zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0);
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0_1[0];
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0_1 = (|_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0);
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h0) == 33'h0));
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2 = (|{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2 = (|_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0);
  assign _zz_WhiteboxerPlugin_logic_csr_access_payload_address = CsrAccessPlugin_logic_fsm_interface_uop;
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h100002040) == 33'h100002000),{((execute_lane1_logic_decoding_decodingBits & 33'h100000044) == 33'h100000004),((execute_lane1_logic_decoding_decodingBits & 33'h100001040) == 33'h100000000)}});
  assign _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100003044) == 33'h100001000));
  assign _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100000010) == 33'h100000000));
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h100000044) == 33'h000000004),{((execute_lane1_logic_decoding_decodingBits & 33'h100002040) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h100001040) == 33'h0)}});
  assign _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100003044) == 33'h000001000));
  assign _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1 = _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2[0];
  assign _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2 = (|_zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1);
  assign _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1[0];
  assign _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1 = (|{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,((execute_lane1_logic_decoding_decodingBits & 33'h000000040) == 33'h0)});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1_1 = (|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane1);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1_1 = (|_zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1);
  assign _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1[0];
  assign _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1 = (|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane1);
  assign _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1 = _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2[0];
  assign _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2 = (|_zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1);
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1[0];
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1 = (|{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1});
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1[0];
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1 = (|_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1);
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h000000010) == 33'h0),{((execute_lane1_logic_decoding_decodingBits & 33'h000002004) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h040000024) == 33'h040000020)}});
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h000000024) == 33'h000000024));
  assign _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1 = _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1[0];
  assign _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1 = 1'b0;
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1_1 = (|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane1);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_1 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_2[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_2 = (|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane1);
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1 = (|_zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1);
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1 = (|_zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1);
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h000002010) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h000005000) == 33'h000001000)});
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2 = (|_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h040000000) == 33'h040000000));
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2 = (|{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1});
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2 = (|_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1);
  assign _zz_WhiteboxerPlugin_logic_loadExecute_data = LsuPlugin_logic_fpwb_payload;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1};
  assign _zz_execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_exponent = execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent;
  assign _zz_execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_exponent = execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent;
  assign _zz_execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent = execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent;
  assign _zz_execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign _zz_BtbPlugin_logic_ras_mem_stack_port = BtbPlugin_logic_ras_write_payload_data;
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[0];
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[1];
  assign _zz_LsuL1Plugin_logic_shared_mem_port = {LsuL1Plugin_logic_shared_write_payload_data_dirty,LsuL1Plugin_logic_shared_write_payload_data_plru_0};
  assign _zz_LsuL1Plugin_logic_writeback_victimBuffer_port = {LsuL1Plugin_logic_writeback_read_slotReadLast_payload_id,LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex};
  assign _zz_PrefetcherRptPlugin_logic_storage_ram_port = {PrefetcherRptPlugin_logic_storage_write_payload_data_missed,{PrefetcherRptPlugin_logic_storage_write_payload_data_advance,{PrefetcherRptPlugin_logic_storage_write_payload_data_score,{PrefetcherRptPlugin_logic_storage_write_payload_data_stride,{PrefetcherRptPlugin_logic_storage_write_payload_data_address,PrefetcherRptPlugin_logic_storage_write_payload_data_tag}}}}};
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[0];
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[1];
  assign _zz_GSharePlugin_logic_mem_banks_0_port = {GSharePlugin_logic_mem_writes_0_payload_data_3,{GSharePlugin_logic_mem_writes_0_payload_data_2,{GSharePlugin_logic_mem_writes_0_payload_data_1,GSharePlugin_logic_mem_writes_0_payload_data_0}}};
  assign _zz_BtbPlugin_logic_mem_port = {{BtbPlugin_logic_memDp_wp_payload_data_1_isPop,{BtbPlugin_logic_memDp_wp_payload_data_1_isPush,{BtbPlugin_logic_memDp_wp_payload_data_1_isBranch,{BtbPlugin_logic_memDp_wp_payload_data_1_pcTarget,{BtbPlugin_logic_memDp_wp_payload_data_1_sliceLow,BtbPlugin_logic_memDp_wp_payload_data_1_hash}}}}},{BtbPlugin_logic_memDp_wp_payload_data_0_isPop,{BtbPlugin_logic_memDp_wp_payload_data_0_isPush,{BtbPlugin_logic_memDp_wp_payload_data_0_isBranch,{BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget,{BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow,BtbPlugin_logic_memDp_wp_payload_data_0_hash}}}}}};
  assign _zz_LsuPlugin_logic_storeBuffer_ops_mem_port_2 = {LsuPlugin_logic_storeBuffer_push_payload_op_storeId,{LsuPlugin_logic_storeBuffer_push_payload_op_size,{LsuPlugin_logic_storeBuffer_push_payload_op_data,LsuPlugin_logic_storeBuffer_push_payload_op_address}}};
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[4 : 3];
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[4 : 3];
  assign _zz_60 = {_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1,_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0};
  assign _zz_62 = {_zz_23[2],{_zz_23[1],_zz_23[0]}};
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[4 : 3];
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[4 : 3];
  assign _zz_64 = {FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH[1],FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH[0]};
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1 = fetch_logic_ctrls_2_down_Fetch_WORD_PC[2 : 1];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28 = AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 10];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30 = {AlignerPlugin_logic_extractors_1_ctx_instruction[12],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]};
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 0];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 1];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_5 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_7 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_67 = {FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[2],{FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[1],FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[0]}};
  assign _zz_DispatchPlugin_logic_candidates_1_age_1 = (DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1);
  assign _zz_DispatchPlugin_logic_candidates_2_age_1 = {(DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1),(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1)};
  assign _zz_DispatchPlugin_logic_slotsFeeds_fit_1 = {(! DispatchPlugin_logic_candidates_2_moving),(! DispatchPlugin_logic_candidates_1_moving)};
  assign _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1 = {DispatchPlugin_logic_candidates_2_ctx_valid,{DispatchPlugin_logic_candidates_1_ctx_valid,DispatchPlugin_logic_candidates_0_ctx_valid}};
  assign _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1 = {decode_ctrls_1_up_LANE_SEL_1,decode_ctrls_1_up_LANE_SEL_0};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[11],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[12],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[13],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[14],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[15],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[16],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[17],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[18],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[19],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[22],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[23],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[24],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[25],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[26],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[27],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[28],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[29],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[30],execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_1 = early0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_2 = early0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_3 = {early0_BarrelShifterPlugin_logic_shift_shifted[11],{early0_BarrelShifterPlugin_logic_shift_shifted[12],{early0_BarrelShifterPlugin_logic_shift_shifted[13],{early0_BarrelShifterPlugin_logic_shift_shifted[14],{early0_BarrelShifterPlugin_logic_shift_shifted[15],{early0_BarrelShifterPlugin_logic_shift_shifted[16],{early0_BarrelShifterPlugin_logic_shift_shifted[17],{early0_BarrelShifterPlugin_logic_shift_shifted[18],{early0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_5,_zz_early0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_4 = early0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_5 = early0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_6 = {early0_BarrelShifterPlugin_logic_shift_shifted[22],{early0_BarrelShifterPlugin_logic_shift_shifted[23],{early0_BarrelShifterPlugin_logic_shift_shifted[24],{early0_BarrelShifterPlugin_logic_shift_shifted[25],{early0_BarrelShifterPlugin_logic_shift_shifted[26],{early0_BarrelShifterPlugin_logic_shift_shifted[27],{early0_BarrelShifterPlugin_logic_shift_shifted[28],{early0_BarrelShifterPlugin_logic_shift_shifted[29],{early0_BarrelShifterPlugin_logic_shift_shifted[30],early0_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[9];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[10];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[11],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[12],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[13],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[14],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[15],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[16],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[17],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[18],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[19],{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_late0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[20];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[21];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[22],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[23],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[24],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[25],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[26],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[27],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[28],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[29],{execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[30],execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_1 = late0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_2 = late0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_3 = {late0_BarrelShifterPlugin_logic_shift_shifted[11],{late0_BarrelShifterPlugin_logic_shift_shifted[12],{late0_BarrelShifterPlugin_logic_shift_shifted[13],{late0_BarrelShifterPlugin_logic_shift_shifted[14],{late0_BarrelShifterPlugin_logic_shift_shifted[15],{late0_BarrelShifterPlugin_logic_shift_shifted[16],{late0_BarrelShifterPlugin_logic_shift_shifted[17],{late0_BarrelShifterPlugin_logic_shift_shifted[18],{late0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_late0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_late0_BarrelShifterPlugin_logic_shift_patched_5,_zz_late0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_4 = late0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_5 = late0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_6 = {late0_BarrelShifterPlugin_logic_shift_shifted[22],{late0_BarrelShifterPlugin_logic_shift_shifted[23],{late0_BarrelShifterPlugin_logic_shift_shifted[24],{late0_BarrelShifterPlugin_logic_shift_shifted[25],{late0_BarrelShifterPlugin_logic_shift_shifted[26],{late0_BarrelShifterPlugin_logic_shift_shifted[27],{late0_BarrelShifterPlugin_logic_shift_shifted[28],{late0_BarrelShifterPlugin_logic_shift_shifted[29],{late0_BarrelShifterPlugin_logic_shift_shifted[30],late0_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[9];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[10];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[11],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[12],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[13],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[14],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[15],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[16],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[17],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[18],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[19],{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early1_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[20];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[21];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[22],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[23],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[24],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[25],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[26],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[27],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[28],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[29],{execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[30],execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_1 = early1_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_2 = early1_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_3 = {early1_BarrelShifterPlugin_logic_shift_shifted[11],{early1_BarrelShifterPlugin_logic_shift_shifted[12],{early1_BarrelShifterPlugin_logic_shift_shifted[13],{early1_BarrelShifterPlugin_logic_shift_shifted[14],{early1_BarrelShifterPlugin_logic_shift_shifted[15],{early1_BarrelShifterPlugin_logic_shift_shifted[16],{early1_BarrelShifterPlugin_logic_shift_shifted[17],{early1_BarrelShifterPlugin_logic_shift_shifted[18],{early1_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early1_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early1_BarrelShifterPlugin_logic_shift_patched_5,_zz_early1_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_4 = early1_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_5 = early1_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_6 = {early1_BarrelShifterPlugin_logic_shift_shifted[22],{early1_BarrelShifterPlugin_logic_shift_shifted[23],{early1_BarrelShifterPlugin_logic_shift_shifted[24],{early1_BarrelShifterPlugin_logic_shift_shifted[25],{early1_BarrelShifterPlugin_logic_shift_shifted[26],{early1_BarrelShifterPlugin_logic_shift_shifted[27],{early1_BarrelShifterPlugin_logic_shift_shifted[28],{early1_BarrelShifterPlugin_logic_shift_shifted[29],{early1_BarrelShifterPlugin_logic_shift_shifted[30],early1_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[9];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[10];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[11],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[12],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[13],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[14],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[15],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[16],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[17],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[18],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[19],{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_5,_zz_late1_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[20];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[21];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[22],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[23],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[24],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[25],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[26],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[27],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[28],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[29],{execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[30],execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_1 = late1_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_2 = late1_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_3 = {late1_BarrelShifterPlugin_logic_shift_shifted[11],{late1_BarrelShifterPlugin_logic_shift_shifted[12],{late1_BarrelShifterPlugin_logic_shift_shifted[13],{late1_BarrelShifterPlugin_logic_shift_shifted[14],{late1_BarrelShifterPlugin_logic_shift_shifted[15],{late1_BarrelShifterPlugin_logic_shift_shifted[16],{late1_BarrelShifterPlugin_logic_shift_shifted[17],{late1_BarrelShifterPlugin_logic_shift_shifted[18],{late1_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_late1_BarrelShifterPlugin_logic_shift_patched_4,{_zz_late1_BarrelShifterPlugin_logic_shift_patched_5,_zz_late1_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_4 = late1_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_5 = late1_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_6 = {late1_BarrelShifterPlugin_logic_shift_shifted[22],{late1_BarrelShifterPlugin_logic_shift_shifted[23],{late1_BarrelShifterPlugin_logic_shift_shifted[24],{late1_BarrelShifterPlugin_logic_shift_shifted[25],{late1_BarrelShifterPlugin_logic_shift_shifted[26],{late1_BarrelShifterPlugin_logic_shift_shifted[27],{late1_BarrelShifterPlugin_logic_shift_shifted[28],{late1_BarrelShifterPlugin_logic_shift_shifted[29],{late1_BarrelShifterPlugin_logic_shift_shifted[30],late1_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts = 1'b1;
  assign _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_1 = fetch_logic_ctrls_0_down_Fetch_WORD_PC[5 : 5];
  assign _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_2 = 1'b0;
  assign _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_3 = fetch_logic_ctrls_0_down_Fetch_WORD_PC[5 : 5];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[7];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[8];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[9],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[10],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[11],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[12],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[13],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[14],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[15],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[16],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[17],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[18];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[19];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[20],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[21],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[22],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[23],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[24],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[25],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[26],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[27],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[28],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[29];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[30];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[31],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[32],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[33],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[34],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[35],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[36],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[37],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[38],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[39],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[40];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[41];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[42],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[43],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[44],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[45],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[46],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[47],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[48],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[49],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[50],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[51];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[52];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[53],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[54],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[55],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[56],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[57],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[58],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[59],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[60],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[61],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[62];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[63];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[64],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[65],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[66],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[67],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[68],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[69],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[70],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[71],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[72],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[73];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[74];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[75],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[76],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[77],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[78],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[79],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[80],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[81],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[82],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[83],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[84];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[85];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[86],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[87],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[88],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[89],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[90],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[91],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[92],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[93],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[94],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26}}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[95];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[96];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26 = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[97],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[98],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[99],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[100],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[101],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[102],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[103],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[104],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[105],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28}}}}}}}}}};
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[106];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28 = FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[107];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_42) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_57) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_59) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_61) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_65) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_1 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_2 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_8) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_11) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_13) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_15) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_19) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_26) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_28) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_30) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_34) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100_2 = (((((FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[1] || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_1) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_3) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_4) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_6);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_43) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_58) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_59) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_62) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_66) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_1 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_2 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_9) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_12) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_13) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_16) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_20) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_27) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_28) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_31) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_35) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101_2 = (((((FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[2] || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_2) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_3) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_5) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_6);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_31) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_37) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_45) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_60) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_61) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_62);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_1 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_2 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_1) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_2) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_3) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_7) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_8) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_9) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_14) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_15) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_16) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_22) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_29) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_30);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102_2 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[4];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_35) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_37) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_49) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_64) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_65) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_66);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_1 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_2 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_4) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_5) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_6) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_7) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_8) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_9) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_18) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_19) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_20) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_22) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_33) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_34);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103_2 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[8];
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_41) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_42) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_43) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_45) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_49) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104_1 = (((((((((((((((FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[16] || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_11) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_12) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_13) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_14) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_15) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_16) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_18) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_19) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_20) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_22) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105 = ((((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_35) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_37) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_41) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_42) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_43) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_45) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_49) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105_1 = (((((((((FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[32] || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_26) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_27) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_28) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_29) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_30) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_31) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_33) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_34);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106 = ((((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106_1 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_66) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_68) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_72) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_73) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_74) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_76) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_80) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83);
  assign _zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106_1 = (((((((((FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[64] || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_57) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_58) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_59) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_60) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_61) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_62) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_64) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_65);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[7];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[8];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2 = {FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[9],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[10],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[11],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[12],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[13],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[14],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[15],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[16],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[17],{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3,{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4,_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5}}}}}}}}}}};
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[18];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[19];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5 = {FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[20],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[21],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[22],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[23],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[24],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[25],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[26],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[27],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[28],{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6,{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7,_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8}}}}}}}}}}};
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[29];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[30];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8 = {FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[31],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[32],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[33],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[34],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[35],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[36],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[37],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[38],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[39],{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9,{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10,_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11}}}}}}}}}}};
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[40];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10 = FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[41];
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11 = {FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[42],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[43],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[44],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[45],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[46],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[47],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[48],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[49],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[50],FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[51]}}}}}}}}};
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123 = (((((((((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[1] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_77) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_78) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_80) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_81) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_83) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_85) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_88) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_90);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124 = (((((((((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[2] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_77) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_79) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_80) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_82) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_83) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_86) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_89) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_90);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125 = (((((((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[4] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_78) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_79) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_80) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_84) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_85) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_86) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126 = (((((((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[8] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_81) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_82) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_83) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_84) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_85) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_86) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127 = ((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[16] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_88) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_89);
  assign _zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128 = ((((_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[32] || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_103) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_104) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_105) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_106);
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask = AlignerPlugin_logic_usedMask_0[4];
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_1 = (! AlignerPlugin_logic_usedMask_0[3]);
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_2 = (AlignerPlugin_logic_scanners_2_valid && (! AlignerPlugin_logic_usedMask_0[2]));
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_3 = (AlignerPlugin_logic_scanners_1_valid && (! AlignerPlugin_logic_usedMask_0[1]));
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_4 = (AlignerPlugin_logic_scanners_0_valid && (! AlignerPlugin_logic_usedMask_0[0]));
  assign _zz_AlignerPlugin_logic_extractors_0_redo_9 = AlignerPlugin_logic_scanners_0_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_10 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_11 = AlignerPlugin_logic_scanners_1_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_12 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_13 = AlignerPlugin_logic_scanners_2_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_14 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_15 = AlignerPlugin_logic_scanners_3_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_16 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_17 = AlignerPlugin_logic_scanners_4_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_18 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_19 = AlignerPlugin_logic_scanners_5_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_20 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_21 = AlignerPlugin_logic_scanners_6_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_22 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_23 = AlignerPlugin_logic_scanners_7_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_24 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask = AlignerPlugin_logic_scanners_0_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_1 = AlignerPlugin_logic_scanners_0_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_2 = AlignerPlugin_logic_scanners_1_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_3 = AlignerPlugin_logic_scanners_1_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_4 = AlignerPlugin_logic_scanners_2_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_5 = AlignerPlugin_logic_scanners_2_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_6 = AlignerPlugin_logic_scanners_3_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_7 = AlignerPlugin_logic_scanners_3_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_8 = AlignerPlugin_logic_scanners_4_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_9 = AlignerPlugin_logic_scanners_4_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_10 = AlignerPlugin_logic_scanners_5_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_11 = AlignerPlugin_logic_scanners_5_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_12 = AlignerPlugin_logic_scanners_6_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_13 = AlignerPlugin_logic_scanners_6_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_14 = AlignerPlugin_logic_scanners_7_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_15 = AlignerPlugin_logic_scanners_7_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask = AlignerPlugin_logic_usedMask_1[4];
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_1 = (! AlignerPlugin_logic_usedMask_1[3]);
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_2 = (AlignerPlugin_logic_scanners_2_valid && (! AlignerPlugin_logic_usedMask_1[2]));
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_3 = (AlignerPlugin_logic_scanners_1_valid && (! AlignerPlugin_logic_usedMask_1[1]));
  assign _zz_AlignerPlugin_logic_extractors_1_redo_8 = AlignerPlugin_logic_scanners_1_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_9 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_10 = AlignerPlugin_logic_scanners_2_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_11 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_12 = AlignerPlugin_logic_scanners_3_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_13 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_14 = AlignerPlugin_logic_scanners_4_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_15 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_16 = AlignerPlugin_logic_scanners_5_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_17 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_18 = AlignerPlugin_logic_scanners_6_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_19 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask = AlignerPlugin_logic_scanners_1_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_1 = AlignerPlugin_logic_scanners_1_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_2 = AlignerPlugin_logic_scanners_2_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_3 = AlignerPlugin_logic_scanners_2_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_4 = AlignerPlugin_logic_scanners_3_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_5 = AlignerPlugin_logic_scanners_3_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_6 = AlignerPlugin_logic_scanners_4_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_7 = AlignerPlugin_logic_scanners_4_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_8 = AlignerPlugin_logic_scanners_5_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_9 = AlignerPlugin_logic_scanners_5_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_10 = AlignerPlugin_logic_scanners_6_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_11 = AlignerPlugin_logic_scanners_6_checker_0_required;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = {_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24 = AlignerPlugin_logic_extractors_0_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = AlignerPlugin_logic_extractors_0_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31 = 7'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32 = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23 = {_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12,AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 3]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24 = AlignerPlugin_logic_extractors_1_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25 = AlignerPlugin_logic_extractors_1_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31 = 7'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32 = AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34 = AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7];
  assign _zz_LsuPlugin_logic_onCtrl_wb_hits = (LsuPlugin_logic_storeBuffer_slots_4_tag == LsuPlugin_logic_onCtrl_wb_tag);
  assign _zz_LsuPlugin_logic_onCtrl_wb_hits_1 = (LsuPlugin_logic_storeBuffer_slots_3_valid && (LsuPlugin_logic_storeBuffer_slots_3_tag == LsuPlugin_logic_onCtrl_wb_tag));
  assign _zz_LsuPlugin_logic_onCtrl_wb_hits_2 = (LsuPlugin_logic_storeBuffer_slots_2_valid && (LsuPlugin_logic_storeBuffer_slots_2_tag == LsuPlugin_logic_onCtrl_wb_tag));
  assign _zz_LsuPlugin_logic_onCtrl_wb_hits_3 = {(LsuPlugin_logic_storeBuffer_slots_1_valid && (LsuPlugin_logic_storeBuffer_slots_1_tag == LsuPlugin_logic_onCtrl_wb_tag)),(LsuPlugin_logic_storeBuffer_slots_0_valid && (LsuPlugin_logic_storeBuffer_slots_0_tag == LsuPlugin_logic_onCtrl_wb_tag))};
  assign _zz_execute_ctrl4_down_LsuL1_ABORD_lane0 = ((! execute_ctrl4_up_LANE_SEL_lane0) || execute_lane0_ctrls_4_upIsCancel);
  assign _zz_execute_ctrl4_down_LsuL1_ABORD_lane0_1 = (! execute_ctrl4_down_LsuL1_FLUSH_lane0);
  assign _zz_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0 = (execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0);
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[0];
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_1 = {FpuPackerPlugin_logic_s0_remapped_0_mantissa,{FpuPackerPlugin_logic_s0_remapped_0_exponent,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_2,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_3}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_4 = 71'h0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_5 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[1];
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_6 = {FpuPackerPlugin_logic_s0_remapped_1_mantissa,{FpuPackerPlugin_logic_s0_remapped_1_exponent,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_7,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_8}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_9 = 71'h0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_10 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[2];
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_11 = {FpuPackerPlugin_logic_s0_remapped_2_mantissa,{FpuPackerPlugin_logic_s0_remapped_2_exponent,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_12,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_13}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_14 = 71'h0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_15 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[3];
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_16 = {FpuPackerPlugin_logic_s0_remapped_3_mantissa,{FpuPackerPlugin_logic_s0_remapped_3_exponent,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_17,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_18}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_19 = 71'h0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_20 = {FpuPackerPlugin_logic_s0_remapped_4_exponent,{FpuPackerPlugin_logic_s0_remapped_4_sign,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_21,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_22}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_23 = {FpuPackerPlugin_logic_s0_remapped_5_exponent,{FpuPackerPlugin_logic_s0_remapped_5_sign,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_24,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_25}}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_2 = FpuPackerPlugin_logic_s0_remapped_0_sign;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_3 = {FpuPackerPlugin_logic_s0_remapped_0_quiet,FpuPackerPlugin_logic_s0_remapped_0_mode};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_7 = FpuPackerPlugin_logic_s0_remapped_1_sign;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_8 = {FpuPackerPlugin_logic_s0_remapped_1_quiet,FpuPackerPlugin_logic_s0_remapped_1_mode};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_12 = FpuPackerPlugin_logic_s0_remapped_2_sign;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_13 = {FpuPackerPlugin_logic_s0_remapped_2_quiet,FpuPackerPlugin_logic_s0_remapped_2_mode};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_17 = FpuPackerPlugin_logic_s0_remapped_3_sign;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_18 = {FpuPackerPlugin_logic_s0_remapped_3_quiet,FpuPackerPlugin_logic_s0_remapped_3_mode};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_21 = FpuPackerPlugin_logic_s0_remapped_4_quiet;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_22 = FpuPackerPlugin_logic_s0_remapped_4_mode;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_24 = FpuPackerPlugin_logic_s0_remapped_5_quiet;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_25 = FpuPackerPlugin_logic_s0_remapped_5_mode;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1 = FpuUnpackerPlugin_logic_packPort_cmd_format;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_1 = 1'b0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_2 = FpuMulPlugin_logic_packPort_cmd_format;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_3 = 1'b0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_4 = FpuSqrtPlugin_logic_packPort_cmd_format;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_5 = 1'b0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_6 = FpuXxPlugin_logic_packPort_cmd_format;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_7 = 1'b0;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX = FpuUnpackerPlugin_logic_packPort_cmd_flags_NV;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_1 = {FpuUnpackerPlugin_logic_packPort_cmd_flags_DZ,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_2,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_3}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_4 = FpuMulPlugin_logic_packPort_cmd_flags_NV;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_5 = {FpuMulPlugin_logic_packPort_cmd_flags_DZ,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_6,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_7}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_8 = FpuSqrtPlugin_logic_packPort_cmd_flags_NV;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_9 = {FpuSqrtPlugin_logic_packPort_cmd_flags_DZ,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_10,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_11}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_12 = FpuXxPlugin_logic_packPort_cmd_flags_NV;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_13 = {FpuXxPlugin_logic_packPort_cmd_flags_DZ,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_14,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_15}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_16 = FpuDivPlugin_logic_packPort_cmd_flags_DZ;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_17 = {FpuDivPlugin_logic_packPort_cmd_flags_OF,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_18,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_19}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_20 = FpuAddSharedPlugin_logic_packPort_cmd_flags_DZ;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_21 = {FpuAddSharedPlugin_logic_packPort_cmd_flags_OF,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_22,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_23}};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_2 = FpuUnpackerPlugin_logic_packPort_cmd_flags_OF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_3 = {FpuUnpackerPlugin_logic_packPort_cmd_flags_UF,FpuUnpackerPlugin_logic_packPort_cmd_flags_NX};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_6 = FpuMulPlugin_logic_packPort_cmd_flags_OF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_7 = {FpuMulPlugin_logic_packPort_cmd_flags_UF,FpuMulPlugin_logic_packPort_cmd_flags_NX};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_10 = FpuSqrtPlugin_logic_packPort_cmd_flags_OF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_11 = {FpuSqrtPlugin_logic_packPort_cmd_flags_UF,FpuSqrtPlugin_logic_packPort_cmd_flags_NX};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_14 = FpuXxPlugin_logic_packPort_cmd_flags_OF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_15 = {FpuXxPlugin_logic_packPort_cmd_flags_UF,FpuXxPlugin_logic_packPort_cmd_flags_NX};
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_18 = FpuDivPlugin_logic_packPort_cmd_flags_UF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_19 = FpuDivPlugin_logic_packPort_cmd_flags_NX;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_22 = FpuAddSharedPlugin_logic_packPort_cmd_flags_UF;
  assign _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_23 = FpuAddSharedPlugin_logic_packPort_cmd_flags_NX;
  assign _zz_execute_lane0_api_hartsInflight = (! execute_ctrl9_down_COMPLETED_lane0);
  assign _zz_execute_lane0_api_hartsInflight_1 = (execute_ctrl8_up_LANE_SEL_lane0 && (! execute_ctrl8_down_COMPLETED_lane0));
  assign _zz_execute_lane0_api_hartsInflight_2 = 1'b1;
  assign _zz_execute_lane0_api_hartsInflight_3 = ((execute_ctrl7_up_LANE_SEL_lane0 && (! execute_ctrl7_down_COMPLETED_lane0)) && 1'b1);
  assign _zz_execute_lane0_api_hartsInflight_4 = ((execute_ctrl6_up_LANE_SEL_lane0 && (! execute_ctrl6_down_COMPLETED_lane0)) && 1'b1);
  assign _zz_execute_lane0_api_hartsInflight_5 = {((execute_ctrl5_up_LANE_SEL_lane0 && (! execute_ctrl5_down_COMPLETED_lane0)) && 1'b1),{(execute_ctrl4_up_LANE_SEL_lane0 && 1'b1),{(execute_ctrl3_up_LANE_SEL_lane0 && _zz_execute_lane0_api_hartsInflight_6),{_zz_execute_lane0_api_hartsInflight_7,_zz_execute_lane0_api_hartsInflight_8}}}};
  assign _zz_execute_lane0_api_hartsInflight_6 = 1'b1;
  assign _zz_execute_lane0_api_hartsInflight_7 = (execute_ctrl2_up_LANE_SEL_lane0 && 1'b1);
  assign _zz_execute_lane0_api_hartsInflight_8 = (execute_ctrl1_up_LANE_SEL_lane0 && 1'b1);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_1 = 32'h00006004;
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00005004);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_3 = 32'h00001000;
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_4 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0_5 = 32'h00002000;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_1 = 32'h00000064;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h08000070);
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_3 = 32'h08000020;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000078) == 32'h00000020);
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_5 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h10000070) == 32'h00000020);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_2 = 32'h00002050;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000070) == 32'h00000030);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006040) == 32'h00004000);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00400028) == 32'h00400000),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000228) == 32'h00000200),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RD_ENABLE_0_6) == 32'h00000004),{(_zz_decode_ctrls_1_down_RD_ENABLE_0_7 == _zz_decode_ctrls_1_down_RD_ENABLE_0_8),{_zz_decode_ctrls_1_down_RD_ENABLE_0_9,{_zz_decode_ctrls_1_down_RD_ENABLE_0_10,_zz_decode_ctrls_1_down_RD_ENABLE_0_11}}}}}};
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_6 = 32'h0000200c;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00800028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_8 = 32'h00800000;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000828) == 32'h00000800);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h000000a8) == 32'h00000080);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h01000028) == 32'h01000000),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000128) == 32'h00000100),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RD_ENABLE_0_12) == 32'h00000400),{(_zz_decode_ctrls_1_down_RD_ENABLE_0_13 == _zz_decode_ctrls_1_down_RD_ENABLE_0_14),(_zz_decode_ctrls_1_down_RD_ENABLE_0_15 == _zz_decode_ctrls_1_down_RD_ENABLE_0_16)}}}};
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_12 = 32'h00000428;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00004028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_14 = 32'h0;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_15 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00100028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_16 = 32'h0;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0 = 32'h0000007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000107f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_2 = 32'h00001073;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000605f) == 32'h00002007),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000705b) == 32'h00002003),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_6) == 32'h00000023),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_7 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_8),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_9,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_10,_zz_decode_ctrls_1_down_Decode_LEGAL_0_11}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_6 = 32'h0000603f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_8 = 32'h00000003;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000506f) == 32'h00000003);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000306f) == 32'h00000003);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000307f) == 32'h00003013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000707b) == 32'h00000063),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_12) == 32'h0000000f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_13 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_14),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_15,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_16,_zz_decode_ctrls_1_down_Decode_LEGAL_0_17}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_12 = 32'h0000607f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000717f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_14 = 32'h00006113;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000787f) == 32'h00006813);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_16 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000727f) == 32'h00006213);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_17 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000747f) == 32'h00006413),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h000070ff) == 32'h00006093),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_18) == 32'h00000053),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_19 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_20),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_21,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_22,_zz_decode_ctrls_1_down_Decode_LEGAL_0_23}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_18 = 32'he400007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_19 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h1800707f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_20 = 32'h0000202f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_21 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc00007f) == 32'h00000033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_22 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'he800707f) == 32'h0800202f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_23 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h7c00607f) == 32'h20000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h7c00507f) == 32'h20000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_24) == 32'h20000053),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_25 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_26),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_27,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_28,_zz_decode_ctrls_1_down_Decode_LEGAL_0_29}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_24 = 32'hf400607f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_25 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc00305f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_26 = 32'h00001013;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_27 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbc00707f) == 32'h00005013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_28 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00005033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_29 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00807fff) == 32'h00806013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h01007fff) == 32'h01006013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_30) == 32'h00406013),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_31 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_32),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_33,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_34,_zz_decode_ctrls_1_down_Decode_LEGAL_0_35}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_30 = 32'h00407fff;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_31 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hede0007f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_32 = 32'hc0000053;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_33 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00000033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_34 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfdf0007f) == 32'h58000053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_35 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h7ff0007f) == 32'h42000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h7ff0007f) == 32'h40100053),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_36) == 32'h00006013),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_37 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_38),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_39,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_40,_zz_decode_ctrls_1_down_Decode_LEGAL_0_41}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_36 = 32'h01c07fff;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_37 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hf9f0707f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_38 = 32'h1000202f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_39 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfdf0707f) == 32'he0001053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_40 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'heff0707f) == 32'he0000053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_41 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffefffff) == 32'h00000073),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffffffff) == 32'h10500073),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffffffff) == 32'h30200073)}};
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1_1 = 32'h00006004;
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00005004);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1_3 = 32'h00001000;
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1_4 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002050);
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_1_5 = 32'h00002000;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1_1 = 32'h00000064;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h08000070);
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1_3 = 32'h08000020;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000078) == 32'h00000020);
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_1_5 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h10000070) == 32'h00000020);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002050);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_2 = 32'h00002050;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000070) == 32'h00000030);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006040) == 32'h00004000);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00400028) == 32'h00400000),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000228) == 32'h00000200),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_RD_ENABLE_1_6) == 32'h00000004),{(_zz_decode_ctrls_1_down_RD_ENABLE_1_7 == _zz_decode_ctrls_1_down_RD_ENABLE_1_8),{_zz_decode_ctrls_1_down_RD_ENABLE_1_9,{_zz_decode_ctrls_1_down_RD_ENABLE_1_10,_zz_decode_ctrls_1_down_RD_ENABLE_1_11}}}}}};
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_6 = 32'h0000200c;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00800028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_8 = 32'h00800000;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000828) == 32'h00000800);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h000000a8) == 32'h00000080);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h01000028) == 32'h01000000),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000128) == 32'h00000100),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_RD_ENABLE_1_12) == 32'h00000400),{(_zz_decode_ctrls_1_down_RD_ENABLE_1_13 == _zz_decode_ctrls_1_down_RD_ENABLE_1_14),(_zz_decode_ctrls_1_down_RD_ENABLE_1_15 == _zz_decode_ctrls_1_down_RD_ENABLE_1_16)}}}};
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_12 = 32'h00000428;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00004028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_14 = 32'h0;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_15 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00100028);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_1_16 = 32'h0;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1 = 32'h0000007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000107f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_2 = 32'h00001073;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000605f) == 32'h00002007),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000705b) == 32'h00002003),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_6) == 32'h00000023),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_7 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_8),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_9,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_10,_zz_decode_ctrls_1_down_Decode_LEGAL_1_11}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_6 = 32'h0000603f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000207f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_8 = 32'h00000003;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000506f) == 32'h00000003);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000306f) == 32'h00000003);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000307f) == 32'h00003013),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000707b) == 32'h00000063),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_12) == 32'h0000000f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_13 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_14),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_15,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_16,_zz_decode_ctrls_1_down_Decode_LEGAL_1_17}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_12 = 32'h0000607f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000717f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_14 = 32'h00006113;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000787f) == 32'h00006813);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_16 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000727f) == 32'h00006213);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_17 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000747f) == 32'h00006413),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h000070ff) == 32'h00006093),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_18) == 32'h00000053),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_19 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_20),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_21,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_22,_zz_decode_ctrls_1_down_Decode_LEGAL_1_23}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_18 = 32'he400007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_19 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h1800707f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_20 = 32'h0000202f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_21 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfc00007f) == 32'h00000033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_22 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'he800707f) == 32'h0800202f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_23 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h7c00607f) == 32'h20000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h7c00507f) == 32'h20000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_24) == 32'h20000053),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_25 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_26),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_27,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_28,_zz_decode_ctrls_1_down_Decode_LEGAL_1_29}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_24 = 32'hf400607f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_25 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfc00305f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_26 = 32'h00001013;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_27 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbc00707f) == 32'h00005013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_28 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbe00707f) == 32'h00005033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_29 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00807fff) == 32'h00806013),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h01007fff) == 32'h01006013),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_30) == 32'h00406013),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_31 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_32),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_33,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_34,_zz_decode_ctrls_1_down_Decode_LEGAL_1_35}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_30 = 32'h00407fff;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_31 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hede0007f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_32 = 32'hc0000053;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_33 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbe00707f) == 32'h00000033);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_34 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfdf0007f) == 32'h58000053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_35 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h7ff0007f) == 32'h42000053),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h7ff0007f) == 32'h40100053),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1_36) == 32'h00006013),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_37 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_38),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_39,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_40,_zz_decode_ctrls_1_down_Decode_LEGAL_1_41}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_36 = 32'h01c07fff;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_37 = (decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hf9f0707f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_38 = 32'h1000202f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_39 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfdf0707f) == 32'he0001053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_40 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'heff0707f) == 32'he0000053);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_1_41 = {((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffefffff) == 32'h00000073),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffffffff) == 32'h10500073),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffffffff) == 32'h30200073)}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1 = (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1) && (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3 = (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5 = (! execute_ctrl2_down_BYPASSED_AT_3_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_6 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_7 = (! execute_ctrl1_down_BYPASSED_AT_2_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_6 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_7 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_8) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_9 = ((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_10 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_11) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_12 = {(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_18,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_21}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_7 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_8 = (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_10 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_11 = (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_13 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_14 = (! execute_ctrl5_down_BYPASSED_AT_6_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_15 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_16 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_17) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_18 = ((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_19 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_20) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_21 = {(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_22 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_23),(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_24 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_25)};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_16 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_17 = (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_19 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_20 = (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_22 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_23 = (! execute_ctrl2_down_BYPASSED_AT_3_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_24 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_25 = (! execute_ctrl1_down_BYPASSED_AT_2_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_6 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_7 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_8) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_9 = ((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_10 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_11) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_12 = {(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_18,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_21}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_7 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_8 = (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_10 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_11 = (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_13 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_14 = (! execute_ctrl5_down_BYPASSED_AT_6_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_15 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_16 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_17) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_18 = ((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_19 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_20) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_21 = {(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_22 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_23),(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_24 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_25)};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_16 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_17 = (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_19 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_20 = (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_22 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_23 = (! execute_ctrl2_down_BYPASSED_AT_3_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_24 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_25 = (! execute_ctrl1_down_BYPASSED_AT_2_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_1 = (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_3 = (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_4 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS)) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_5 = (! execute_ctrl7_down_BYPASSED_AT_8_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_6 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_7 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_8) && (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID)) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_9 = ((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_10 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_11) && (! execute_ctrl5_down_BYPASSED_AT_6_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_12 = {(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_16,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_19}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_7 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_8 = (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_10 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_11 = (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_13 = (((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS)) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_14 = (! execute_ctrl4_down_BYPASSED_AT_5_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_15 = ((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS)) && (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID)) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_16 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_17 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_18) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_19 = (((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_20 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_21) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_17 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_18 = (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_20 = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_21 = (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_6 = (((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_7 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_8) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_9 = ((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_10 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_11) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_12 = {(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_16,_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_19}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_7 = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_8 = (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_10 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_11 = (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_13 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_14 = (! execute_ctrl5_down_BYPASSED_AT_6_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_15 = ((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_16 = (((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_17 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_18) && (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_19 = {((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_20 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_21) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_22 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_23) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_17 = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_18 = (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_20 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_21 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_22 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_23 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_6 = (((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_7 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_8) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_9 = ((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_10 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_11) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_12 = {(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_16,_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_19}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_7 = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_8 = (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_10 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_11 = (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_13 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_14 = (! execute_ctrl5_down_BYPASSED_AT_6_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_15 = ((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_16 = (((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_17 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_18) && (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_19 = {((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_20 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_21) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_22 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_23) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_17 = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_18 = (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_20 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_21 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_22 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_23 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_1 = (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_3 = (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_4 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_5 = (! execute_ctrl6_down_BYPASSED_AT_7_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_6 = ((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID)) && (! execute_ctrl5_down_BYPASSED_AT_6_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_7 = (((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_8 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_9) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_10 = {((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_11 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_12) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_14),(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_15 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_16)}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_8 = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_9 = (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_11 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_12 = (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_13 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_14 = (! execute_ctrl2_down_BYPASSED_AT_3_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_15 = (((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_16 = (! execute_ctrl1_down_BYPASSED_AT_2_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3 = (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5 = (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_6 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_7 = (((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_8 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_9) && (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_10 = {((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_11 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_12) && (! execute_ctrl5_down_BYPASSED_AT_6_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_16,_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_17}}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_8 = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_9 = (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_11 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_12 = (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_13 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_14 = (! execute_ctrl4_down_BYPASSED_AT_5_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_15 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_16 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_17 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1 = (execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3 = (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5 = (! execute_ctrl8_down_BYPASSED_AT_9_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_6 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_7 = (((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_8 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_9) && (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl6_down_BYPASSED_AT_7_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_10 = {((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_11 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_12) && (! execute_ctrl5_down_BYPASSED_AT_6_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_14),{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_15,{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_16,_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_17}}}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_8 = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_9 = (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_11 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_12 = (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_13 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_14 = (! execute_ctrl4_down_BYPASSED_AT_5_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_15 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_16 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_17 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl8_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_1 = (execute_ctrl8_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_3 = (execute_ctrl7_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_4 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (execute_ctrl6_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_5 = (! execute_ctrl6_down_BYPASSED_AT_7_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_6 = ((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (execute_ctrl5_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID)) && (! execute_ctrl5_down_BYPASSED_AT_6_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_7 = (((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_8 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_9) && (execute_ctrl4_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID)) && (! execute_ctrl4_down_BYPASSED_AT_5_lane0));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_10 = {((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_11 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_12) && (! execute_ctrl3_down_BYPASSED_AT_4_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_13 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_14),(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_15 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_16)}};
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_8 = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl4_up_RD_ENABLE_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_9 = (execute_ctrl4_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_11 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_12 = (execute_ctrl3_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_13 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (execute_ctrl2_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_14 = (! execute_ctrl2_down_BYPASSED_AT_3_lane0);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_15 = (((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (execute_ctrl1_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_16 = (! execute_ctrl1_down_BYPASSED_AT_2_lane0);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_3 = 32'hffd02050;
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_4 = 32'hffd01050;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_4 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1}}};
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_2 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_3 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1}}}};
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_18 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_19 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1}}}};
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_3 = 32'hffd02050;
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_4 = 32'hffd01050;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_4 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1}}};
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_2 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_3 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1}}}};
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_18 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_19 = {_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3,{_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,_zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1}}}};
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_1 = {fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash};
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_2 = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_3 = {fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash};
  assign _zz_AlignerPlugin_logic_buffer_flushIt = 1'b1;
  assign _zz_AlignerPlugin_logic_buffer_flushIt_1 = (early0_EnvPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_AlignerPlugin_logic_buffer_flushIt_2 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_AlignerPlugin_logic_buffer_flushIt_3 = {(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)};
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[0];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[1];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[3];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[4];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[6];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[7];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16 = 32'h0;
  assign _zz_DispatchPlugin_logic_candidates_0_cancel = 1'b1;
  assign _zz_DispatchPlugin_logic_candidates_0_cancel_1 = 1'b1;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4 = DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14 = DispatchPlugin_logic_candidates_1_ctx_valid;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15 = DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_29 = DispatchPlugin_logic_candidates_2_ctx_valid;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2 = DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID,{DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE,{DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17 = DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID,{DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE,{DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4 = DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5 = {DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID,{DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE,{DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID,{DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19 = DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20 = {DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID,{DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE,{DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID,{DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_22}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6 = DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7 = {DispatchPlugin_logic_candidates_1_ctx_hm_TRAP,{DispatchPlugin_logic_candidates_1_ctx_hm_PC,{DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4,{DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3,{DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21 = DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_22 = {DispatchPlugin_logic_candidates_2_ctx_hm_TRAP,{DispatchPlugin_logic_candidates_2_ctx_hm_PC,{DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4,{DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3,{DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_23,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_24}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8 = DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9 = {DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9,{DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5,{DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5,{DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6,{DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_23 = DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_24 = {DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9,{DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5,{DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5,{DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6,{DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_25,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_26}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10 = DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_25 = DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_26 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_27,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_28}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12 = {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13 = {DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC,DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_27 = {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_28 = {DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC,DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED}}};
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1 = {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0};
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3 = {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0};
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4 = DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5 = DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt = 1'b1;
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_3 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt = 1'b1;
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_3 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt = 1'b0;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_1 = (DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge == 1'b0);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_2 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_3 = (DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge < 1'b0);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_4 = ((DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge == 1'b0) && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_5 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_6 = (early1_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_7 = (late0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_8 = {(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}};
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_1 = (DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge == _zz_decode_logic_flushes_1_onLanes_1_doIt);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_2 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_3 = (late0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_4 = (early0_EnvPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_5 = {(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception};
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_6 = TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_7 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_8 = late0_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_9 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_10 = late1_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_11 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_12 = early0_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_13 = 32'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented = COMB_CSR_834;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1 = {COMB_CSR_768,{COMB_CSR_769,{COMB_CSR_3860,{COMB_CSR_3859,{COMB_CSR_3858,{COMB_CSR_3857,{COMB_CSR_1954,{COMB_CSR_1953,{COMB_CSR_1952,COMB_CSR_2047}}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = 32'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = 32'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = 32'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_769) ? 32'h4000112d : 32'h0);
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1 = _zz_execute_ctrl1_down_integer_RS1_lane0[0];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_1 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_2 = _zz_execute_ctrl1_down_integer_RS1_lane0[1];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_3 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_4 = _zz_execute_ctrl1_down_integer_RS1_lane0[2];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_5 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_6 = _zz_execute_ctrl1_down_integer_RS1_lane0[3];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_7 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_8 = _zz_execute_ctrl1_down_integer_RS1_lane0[4];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_9 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_10 = _zz_execute_ctrl1_down_integer_RS1_lane0[5];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_11 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_12 = _zz_execute_ctrl1_down_integer_RS1_lane0[6];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_13 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_14 = _zz_execute_ctrl1_down_integer_RS1_lane0[7];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_15 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1 = _zz_execute_ctrl1_down_integer_RS2_lane0[0];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_1 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_2 = _zz_execute_ctrl1_down_integer_RS2_lane0[1];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_3 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_4 = _zz_execute_ctrl1_down_integer_RS2_lane0[2];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_5 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_6 = _zz_execute_ctrl1_down_integer_RS2_lane0[3];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_7 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_8 = _zz_execute_ctrl1_down_integer_RS2_lane0[4];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_9 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_10 = _zz_execute_ctrl1_down_integer_RS2_lane0[5];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_11 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_12 = _zz_execute_ctrl1_down_integer_RS2_lane0[6];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_13 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_14 = _zz_execute_ctrl1_down_integer_RS2_lane0[7];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_15 = 32'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0 = execute_lane0_bypasser_float_RS1_sel[0];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_1 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_2 = execute_lane0_bypasser_float_RS1_sel[1];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_3 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_4 = execute_lane0_bypasser_float_RS1_sel[2];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_5 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_6 = execute_lane0_bypasser_float_RS1_sel[3];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_7 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_8 = execute_lane0_bypasser_float_RS1_sel[4];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_9 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_10 = execute_lane0_bypasser_float_RS1_sel[5];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_11 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_12 = execute_lane0_bypasser_float_RS1_sel[6];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_13 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS1_lane0_14 = execute_lane0_bypasser_float_RS1_sel[7];
  assign _zz_execute_ctrl1_down_float_RS1_lane0_15 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0 = execute_lane0_bypasser_float_RS2_sel[0];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_1 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_2 = execute_lane0_bypasser_float_RS2_sel[1];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_3 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_4 = execute_lane0_bypasser_float_RS2_sel[2];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_5 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_6 = execute_lane0_bypasser_float_RS2_sel[3];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_7 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_8 = execute_lane0_bypasser_float_RS2_sel[4];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_9 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_10 = execute_lane0_bypasser_float_RS2_sel[5];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_11 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_12 = execute_lane0_bypasser_float_RS2_sel[6];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_13 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS2_lane0_14 = execute_lane0_bypasser_float_RS2_sel[7];
  assign _zz_execute_ctrl1_down_float_RS2_lane0_15 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0 = execute_lane0_bypasser_float_RS3_sel[0];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_1 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_2 = execute_lane0_bypasser_float_RS3_sel[1];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_3 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_4 = execute_lane0_bypasser_float_RS3_sel[2];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_5 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_6 = execute_lane0_bypasser_float_RS3_sel[3];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_7 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_8 = execute_lane0_bypasser_float_RS3_sel[4];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_9 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_10 = execute_lane0_bypasser_float_RS3_sel[5];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_11 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_12 = execute_lane0_bypasser_float_RS3_sel[6];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_13 = 64'h0;
  assign _zz_execute_ctrl1_down_float_RS3_lane0_14 = execute_lane0_bypasser_float_RS3_sel[7];
  assign _zz_execute_ctrl1_down_float_RS3_lane0_15 = 64'h0;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_2 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_3;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_3 = {_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_1,{((execute_lane0_logic_decoding_decodingBits & 33'h100006070) == 33'h100002010),{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h102001070) == 33'h100000030),((execute_lane0_logic_decoding_decodingBits & 33'h100003070) == 33'h100000010)}}}}};
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3 = 33'h000002030;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4 = (execute_lane0_logic_decoding_decodingBits & 33'h000000070);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5 = 33'h000000030;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002024) == 33'h000000024);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_7 = ((execute_lane0_logic_decoding_decodingBits & 33'h000006040) == 33'h000004000);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_8 = {((execute_lane0_logic_decoding_decodingBits & 33'h090000050) == 33'h080000050),{((execute_lane0_logic_decoding_decodingBits & 33'h0000000e4) == 33'h000000080),{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_9) == 33'h000000800),{(_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_10 == _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_11),{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_12,{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_13,_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_14}}}}}};
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_9 = 33'h000000864;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_10 = (execute_lane0_logic_decoding_decodingBits & 33'h000000164);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_11 = 33'h000000100;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_12 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000264) == 33'h000000200);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_13 = ((execute_lane0_logic_decoding_decodingBits & 33'h001000064) == 33'h001000000);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_14 = {((execute_lane0_logic_decoding_decodingBits & 33'h000001064) == 33'h000001000),{((execute_lane0_logic_decoding_decodingBits & 33'h000400064) == 33'h000400000),{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_15) == 33'h000800000),{(_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_16 == _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_17),{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_18,_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_19}}}}};
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_15 = 33'h000800064;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_16 = (execute_lane0_logic_decoding_decodingBits & 33'h000000464);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_17 = 33'h000000400;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_18 = ((execute_lane0_logic_decoding_decodingBits & 33'h000004064) == 33'h0);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_19 = ((execute_lane0_logic_decoding_decodingBits & 33'h000100064) == 33'h0);
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_2 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_6;
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_3 = {_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_5,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0}}}}};
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_18 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_6;
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_19 = {_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_5,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0}}}}};
  assign _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1 = 33'h042000000;
  assign _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_1 = 33'h0d2000010;
  assign _zz_when_ExecuteLanePlugin_l306_2 = (early1_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l306_2_1 = (early0_EnvPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_when_ExecuteLanePlugin_l306_2_2 = ((early0_EnvPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane0) || ((early0_EnvPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane0) && early0_EnvPlugin_logic_flushPort_payload_self));
  assign _zz_when_ExecuteLanePlugin_l306_2_3 = ((CsrAccessPlugin_logic_flushPort_valid && 1'b1) && ((CsrAccessPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane0) || ((CsrAccessPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane0) && CsrAccessPlugin_logic_flushPort_payload_self)));
  assign _zz_when_ExecuteLanePlugin_l306_2_4 = ((early0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early0_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane0) || ((early0_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane0) && early0_BranchPlugin_logic_flushPort_payload_self)));
  assign _zz_when_ExecuteLanePlugin_l306_2_5 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_when_ExecuteLanePlugin_l306_4 = (late0_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l306_4_1 = (LsuPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane0);
  assign _zz_fetch_logic_flushes_0_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_0_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_0_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_0_doIt_3 = {(LsuPlugin_logic_flushPort_valid && 1'b1),((BtbPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && BtbPlugin_logic_flushPort_payload_self)))};
  assign _zz_fetch_logic_flushes_1_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_1_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_1_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_1_doIt_3 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1 = _zz_execute_ctrl1_down_integer_RS1_lane1[0];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_1 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_2 = _zz_execute_ctrl1_down_integer_RS1_lane1[1];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_3 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_4 = _zz_execute_ctrl1_down_integer_RS1_lane1[2];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_5 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_6 = _zz_execute_ctrl1_down_integer_RS1_lane1[3];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_7 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_8 = _zz_execute_ctrl1_down_integer_RS1_lane1[4];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_9 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_10 = _zz_execute_ctrl1_down_integer_RS1_lane1[5];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_11 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_12 = _zz_execute_ctrl1_down_integer_RS1_lane1[6];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_13 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_14 = _zz_execute_ctrl1_down_integer_RS1_lane1[7];
  assign _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_15 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1 = _zz_execute_ctrl1_down_integer_RS2_lane1[0];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_1 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_2 = _zz_execute_ctrl1_down_integer_RS2_lane1[1];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_3 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_4 = _zz_execute_ctrl1_down_integer_RS2_lane1[2];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_5 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_6 = _zz_execute_ctrl1_down_integer_RS2_lane1[3];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_7 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_8 = _zz_execute_ctrl1_down_integer_RS2_lane1[4];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_9 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_10 = _zz_execute_ctrl1_down_integer_RS2_lane1[5];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_11 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_12 = _zz_execute_ctrl1_down_integer_RS2_lane1[6];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_13 = 32'h0;
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_14 = _zz_execute_ctrl1_down_integer_RS2_lane1[7];
  assign _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_15 = 32'h0;
  assign _zz_when_ExecuteLanePlugin_l306_7 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l306_7_1 = (early0_EnvPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l306_7_2 = ((early0_EnvPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane1) && early0_EnvPlugin_logic_flushPort_payload_self);
  assign _zz_when_ExecuteLanePlugin_l306_7_3 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_when_ExecuteLanePlugin_l306_7_4 = ((CsrAccessPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane1) || ((CsrAccessPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane1) && CsrAccessPlugin_logic_flushPort_payload_self));
  assign _zz_when_ExecuteLanePlugin_l306_7_5 = ((early0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early0_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane1) || ((early0_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane1) && early0_BranchPlugin_logic_flushPort_payload_self)));
  assign _zz_when_ExecuteLanePlugin_l306_7_6 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_when_ExecuteLanePlugin_l306_9 = (late0_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l306_9_1 = (LsuPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane1);
  assign _zz_TrapPlugin_logic_initHold = 1'b0;
  assign _zz_TrapPlugin_logic_initHold_1 = 1'b0;
  assign _zz_TrapPlugin_logic_initHold_2 = 1'b0;
  assign BtbPlugin_logic_ras_mem_stack_spinal_port0 = BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_ptr_pop_aheadValue];
  always @(posedge clk) begin
    if(_zz_3) begin
      BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_write_payload_address] <= _zz_BtbPlugin_logic_ras_mem_stack_port;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_0_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_0_memsymbol_read_31, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_30, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_29, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_28, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_27, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_26, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_25, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_24, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_23, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_22, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_21, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_20, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_19, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_18, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_17, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_16, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_15, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_14, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_13, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_12, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_11, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_10, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_9, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_8, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read};
  end
  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[0] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[1] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[2] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[3] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[4] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[5] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[6] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[7] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[63 : 56];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[8] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol8[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[71 : 64];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[9] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol9[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[79 : 72];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[10] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol10[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[87 : 80];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[11] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol11[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[95 : 88];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[12] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol12[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[103 : 96];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[13] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol13[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[111 : 104];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[14] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol14[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[119 : 112];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[15] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol15[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[127 : 120];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[16] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol16[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[135 : 128];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[17] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol17[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[143 : 136];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[18] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol18[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[151 : 144];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[19] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol19[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[159 : 152];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[20] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol20[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[167 : 160];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[21] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol21[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[175 : 168];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[22] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol22[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[183 : 176];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[23] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol23[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[191 : 184];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[24] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol24[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[199 : 192];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[25] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol25[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[207 : 200];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[26] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol26[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[215 : 208];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[27] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol27[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[223 : 216];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[28] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol28[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[231 : 224];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[29] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol29[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[239 : 232];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[30] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol30[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[247 : 240];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[31] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol31[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[255 : 248];
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_0_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read <= LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1 <= LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2 <= LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3 <= LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4 <= LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5 <= LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6 <= LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7 <= LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_8 <= LsuL1Plugin_logic_banks_0_mem_symbol8[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_9 <= LsuL1Plugin_logic_banks_0_mem_symbol9[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_10 <= LsuL1Plugin_logic_banks_0_mem_symbol10[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_11 <= LsuL1Plugin_logic_banks_0_mem_symbol11[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_12 <= LsuL1Plugin_logic_banks_0_mem_symbol12[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_13 <= LsuL1Plugin_logic_banks_0_mem_symbol13[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_14 <= LsuL1Plugin_logic_banks_0_mem_symbol14[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_15 <= LsuL1Plugin_logic_banks_0_mem_symbol15[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_16 <= LsuL1Plugin_logic_banks_0_mem_symbol16[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_17 <= LsuL1Plugin_logic_banks_0_mem_symbol17[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_18 <= LsuL1Plugin_logic_banks_0_mem_symbol18[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_19 <= LsuL1Plugin_logic_banks_0_mem_symbol19[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_20 <= LsuL1Plugin_logic_banks_0_mem_symbol20[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_21 <= LsuL1Plugin_logic_banks_0_mem_symbol21[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_22 <= LsuL1Plugin_logic_banks_0_mem_symbol22[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_23 <= LsuL1Plugin_logic_banks_0_mem_symbol23[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_24 <= LsuL1Plugin_logic_banks_0_mem_symbol24[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_25 <= LsuL1Plugin_logic_banks_0_mem_symbol25[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_26 <= LsuL1Plugin_logic_banks_0_mem_symbol26[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_27 <= LsuL1Plugin_logic_banks_0_mem_symbol27[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_28 <= LsuL1Plugin_logic_banks_0_mem_symbol28[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_29 <= LsuL1Plugin_logic_banks_0_mem_symbol29[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_30 <= LsuL1Plugin_logic_banks_0_mem_symbol30[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_31 <= LsuL1Plugin_logic_banks_0_mem_symbol31[LsuL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_1_memsymbol_read_31, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_30, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_29, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_28, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_27, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_26, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_25, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_24, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_23, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_22, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_21, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_20, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_19, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_18, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_17, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_16, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_15, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_14, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_13, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_12, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_11, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_10, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_9, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_8, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read};
  end
  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[0] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[1] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[2] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[3] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[4] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[5] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[6] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[7] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[63 : 56];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[8] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol8[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[71 : 64];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[9] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol9[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[79 : 72];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[10] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol10[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[87 : 80];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[11] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol11[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[95 : 88];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[12] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol12[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[103 : 96];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[13] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol13[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[111 : 104];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[14] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol14[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[119 : 112];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[15] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol15[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[127 : 120];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[16] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol16[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[135 : 128];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[17] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol17[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[143 : 136];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[18] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol18[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[151 : 144];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[19] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol19[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[159 : 152];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[20] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol20[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[167 : 160];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[21] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol21[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[175 : 168];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[22] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol22[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[183 : 176];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[23] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol23[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[191 : 184];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[24] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol24[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[199 : 192];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[25] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol25[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[207 : 200];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[26] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol26[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[215 : 208];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[27] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol27[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[223 : 216];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[28] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol28[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[231 : 224];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[29] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol29[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[239 : 232];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[30] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol30[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[247 : 240];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[31] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol31[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[255 : 248];
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_banks_1_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read <= LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1 <= LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2 <= LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3 <= LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4 <= LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5 <= LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6 <= LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7 <= LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_8 <= LsuL1Plugin_logic_banks_1_mem_symbol8[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_9 <= LsuL1Plugin_logic_banks_1_mem_symbol9[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_10 <= LsuL1Plugin_logic_banks_1_mem_symbol10[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_11 <= LsuL1Plugin_logic_banks_1_mem_symbol11[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_12 <= LsuL1Plugin_logic_banks_1_mem_symbol12[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_13 <= LsuL1Plugin_logic_banks_1_mem_symbol13[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_14 <= LsuL1Plugin_logic_banks_1_mem_symbol14[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_15 <= LsuL1Plugin_logic_banks_1_mem_symbol15[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_16 <= LsuL1Plugin_logic_banks_1_mem_symbol16[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_17 <= LsuL1Plugin_logic_banks_1_mem_symbol17[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_18 <= LsuL1Plugin_logic_banks_1_mem_symbol18[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_19 <= LsuL1Plugin_logic_banks_1_mem_symbol19[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_20 <= LsuL1Plugin_logic_banks_1_mem_symbol20[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_21 <= LsuL1Plugin_logic_banks_1_mem_symbol21[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_22 <= LsuL1Plugin_logic_banks_1_mem_symbol22[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_23 <= LsuL1Plugin_logic_banks_1_mem_symbol23[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_24 <= LsuL1Plugin_logic_banks_1_mem_symbol24[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_25 <= LsuL1Plugin_logic_banks_1_mem_symbol25[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_26 <= LsuL1Plugin_logic_banks_1_mem_symbol26[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_27 <= LsuL1Plugin_logic_banks_1_mem_symbol27[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_28 <= LsuL1Plugin_logic_banks_1_mem_symbol28[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_29 <= LsuL1Plugin_logic_banks_1_mem_symbol29[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_30 <= LsuL1Plugin_logic_banks_1_mem_symbol30[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_31 <= LsuL1Plugin_logic_banks_1_mem_symbol31[LsuL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_LsuL1Plugin_logic_ways_0_mem_port_1) begin
      LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_0_mem_spinal_port1 <= LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_LsuL1Plugin_logic_ways_1_mem_port_1) begin
      LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_1_mem_spinal_port1 <= LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_10) begin
      LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_write_payload_address] <= _zz_LsuL1Plugin_logic_shared_mem_port;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_shared_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_shared_mem_spinal_port1 <= LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_9) begin
      LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_victimBuffer_port] <= LsuL1Plugin_logic_writeback_read_readedData;
    end
  end

  always @(posedge clk) begin
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1 <= LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_write_word];
    end
  end

  always @(posedge clk) begin
    if(PrefetcherRptPlugin_logic_storage_read_cmd_valid) begin
      PrefetcherRptPlugin_logic_storage_ram_spinal_port0 <= PrefetcherRptPlugin_logic_storage_ram[PrefetcherRptPlugin_logic_storage_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_8) begin
      PrefetcherRptPlugin_logic_storage_ram[PrefetcherRptPlugin_logic_storage_write_payload_address] <= _zz_PrefetcherRptPlugin_logic_storage_ram_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_7) begin
      FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_write_payload_address] <= FetchL1Plugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_banks_0_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_0_mem_spinal_port1 <= FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_6) begin
      FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_write_payload_address] <= FetchL1Plugin_logic_banks_1_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_banks_1_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_1_mem_spinal_port1 <= FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_ways_0_mem_port_1) begin
      FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_ways_0_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_0_mem_spinal_port1 <= FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_ways_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchL1Plugin_logic_ways_1_mem_port_1) begin
      FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_ways_1_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_1_mem_spinal_port1 <= FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_ways_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_5) begin
      FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_write_payload_address] <= FetchL1Plugin_logic_plru_write_payload_data_0;
    end
  end

  always @(posedge clk) begin
    if(FetchL1Plugin_logic_plru_read_cmd_valid) begin
      FetchL1Plugin_logic_plru_mem_spinal_port1 <= FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_4) begin
      GSharePlugin_logic_mem_banks_0[GSharePlugin_logic_mem_writes_0_payload_address] <= _zz_GSharePlugin_logic_mem_banks_0_port;
    end
  end

  always @(posedge clk) begin
    if(fetch_logic_ctrls_0_down_isReady) begin
      GSharePlugin_logic_mem_banks_0_spinal_port1 <= GSharePlugin_logic_mem_banks_0[_zz_GSharePlugin_logic_readRsp_readed_0_0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_mem_spinal_port1 = {_zz_BtbPlugin_logic_memsymbol_read_1, _zz_BtbPlugin_logic_memsymbol_read};
  end
  always @(posedge clk) begin
    if(BtbPlugin_logic_memDp_wp_payload_mask[0] && BtbPlugin_logic_memDp_wp_valid) begin
      BtbPlugin_logic_mem_symbol0[BtbPlugin_logic_memDp_wp_payload_address] <= _zz_BtbPlugin_logic_mem_port[46 : 0];
    end
    if(BtbPlugin_logic_memDp_wp_payload_mask[1] && BtbPlugin_logic_memDp_wp_valid) begin
      BtbPlugin_logic_mem_symbol1[BtbPlugin_logic_memDp_wp_payload_address] <= _zz_BtbPlugin_logic_mem_port[93 : 47];
    end
  end

  always @(posedge clk) begin
    if(BtbPlugin_logic_memDp_rp_cmd_valid) begin
      _zz_BtbPlugin_logic_memsymbol_read <= BtbPlugin_logic_mem_symbol0[BtbPlugin_logic_memDp_rp_cmd_payload];
      _zz_BtbPlugin_logic_memsymbol_read_1 <= BtbPlugin_logic_mem_symbol1[BtbPlugin_logic_memDp_rp_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(LsuPlugin_logic_storeBuffer_ops_pip_node_0_isFiring) begin
      LsuPlugin_logic_storeBuffer_ops_mem_spinal_port0 <= LsuPlugin_logic_storeBuffer_ops_mem[_zz__zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      LsuPlugin_logic_storeBuffer_ops_mem[_zz_LsuPlugin_logic_storeBuffer_ops_mem_port_1] <= _zz_LsuPlugin_logic_storeBuffer_ops_mem_port_2;
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  always @(posedge clk) begin
    if(CsrRamPlugin_logic_readLogic_port_cmd_valid) begin
      CsrRamPlugin_logic_mem_spinal_port1 <= CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_cmd_payload];
    end
  end

  StreamFifo PrefetcherRptPlugin_logic_order_fifo (
    .io_push_valid           (PrefetcherRptPlugin_logic_order_valid                            ), //i
    .io_push_ready           (PrefetcherRptPlugin_logic_order_fifo_io_push_ready               ), //o
    .io_push_payload_address (PrefetcherRptPlugin_logic_order_payload_address[31:0]            ), //i
    .io_push_payload_unique  (PrefetcherRptPlugin_logic_order_payload_unique                   ), //i
    .io_push_payload_from    (PrefetcherRptPlugin_logic_order_payload_from[2:0]                ), //i
    .io_push_payload_to      (PrefetcherRptPlugin_logic_order_payload_to[2:0]                  ), //i
    .io_push_payload_stride  (PrefetcherRptPlugin_logic_order_payload_stride[11:0]             ), //i
    .io_pop_valid            (PrefetcherRptPlugin_logic_order_fifo_io_pop_valid                ), //o
    .io_pop_ready            (PrefetcherRptPlugin_logic_queued_ready                           ), //i
    .io_pop_payload_address  (PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_address[31:0]), //o
    .io_pop_payload_unique   (PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_unique       ), //o
    .io_pop_payload_from     (PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_from[2:0]    ), //o
    .io_pop_payload_to       (PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_to[2:0]      ), //o
    .io_pop_payload_stride   (PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_stride[11:0] ), //o
    .io_flush                (1'b0                                                             ), //i
    .io_occupancy            (PrefetcherRptPlugin_logic_order_fifo_io_occupancy[2:0]           ), //o
    .io_availability         (PrefetcherRptPlugin_logic_order_fifo_io_availability[2:0]        ), //o
    .clk                     (clk                                                              ), //i
    .reset                   (reset                                                            )  //i
  );
  StreamArbiter LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter (
    .io_inputs_0_valid                    (LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_valid                                   ), //i
    .io_inputs_0_ready                    (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_0_ready                       ), //o
    .io_inputs_0_payload_last             (LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_last                            ), //i
    .io_inputs_0_payload_fragment_write   (LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_write                  ), //i
    .io_inputs_0_payload_fragment_id      (LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_id                     ), //i
    .io_inputs_0_payload_fragment_address (LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_address[31:0]          ), //i
    .io_inputs_1_valid                    (LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_valid                                  ), //i
    .io_inputs_1_ready                    (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_1_ready                       ), //o
    .io_inputs_1_payload_last             (LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_last                           ), //i
    .io_inputs_1_payload_fragment_write   (LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_write                 ), //i
    .io_inputs_1_payload_fragment_id      (LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_id                    ), //i
    .io_inputs_1_payload_fragment_address (LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_address[31:0]         ), //i
    .io_output_valid                      (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_valid                         ), //o
    .io_output_ready                      (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_ready                         ), //i
    .io_output_payload_last               (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_last                  ), //o
    .io_output_payload_fragment_write     (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_write        ), //o
    .io_output_payload_fragment_id        (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_id           ), //o
    .io_output_payload_fragment_address   (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_address[31:0]), //o
    .io_chosen                            (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_chosen                               ), //o
    .io_chosenOH                          (LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_chosenOH[1:0]                        ), //o
    .clk                                  (clk                                                                                      ), //i
    .reset                                (reset                                                                                    )  //i
  );
  StreamArbiter_1 FpuUnpackerPlugin_logic_unpacker_arbiter (
    .io_inputs_0_valid        (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid             ), //i
    .io_inputs_0_ready        (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_ready             ), //o
    .io_inputs_0_payload_data (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data[51:0]), //i
    .io_inputs_1_valid        (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_valid             ), //i
    .io_inputs_1_ready        (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_ready             ), //o
    .io_inputs_1_payload_data (FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_payload_data[51:0]), //i
    .io_output_valid          (FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_valid               ), //o
    .io_output_ready          (1'b1                                                                   ), //i
    .io_output_payload_data   (FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_payload_data[51:0]  ), //o
    .io_chosen                (FpuUnpackerPlugin_logic_unpacker_arbiter_io_chosen                     ), //o
    .io_chosenOH              (FpuUnpackerPlugin_logic_unpacker_arbiter_io_chosenOH[1:0]              ), //o
    .clk                      (clk                                                                    ), //i
    .reset                    (reset                                                                  )  //i
  );
  DivRadix early0_DivPlugin_logic_processing_div (
    .io_flush                  (execute_ctrl2_down_isReady                                          ), //i
    .io_cmd_valid              (early0_DivPlugin_logic_processing_div_io_cmd_valid                  ), //i
    .io_cmd_ready              (early0_DivPlugin_logic_processing_div_io_cmd_ready                  ), //o
    .io_cmd_payload_a          (early0_DivPlugin_logic_processing_a[63:0]                           ), //i
    .io_cmd_payload_b          (early0_DivPlugin_logic_processing_b[63:0]                           ), //i
    .io_cmd_payload_normalized (early0_DivPlugin_logic_processing_div_io_cmd_payload_normalized     ), //i
    .io_cmd_payload_iterations (early0_DivPlugin_logic_processing_div_io_cmd_payload_iterations[4:0]), //i
    .io_rsp_valid              (early0_DivPlugin_logic_processing_div_io_rsp_valid                  ), //o
    .io_rsp_ready              (1'b0                                                                ), //i
    .io_rsp_payload_result     (early0_DivPlugin_logic_processing_div_io_rsp_payload_result[63:0]   ), //o
    .io_rsp_payload_remain     (early0_DivPlugin_logic_processing_div_io_rsp_payload_remain[63:0]   ), //o
    .clk                       (clk                                                                 ), //i
    .reset                     (reset                                                               )  //i
  );
  StreamArbiter_2 LsuPlugin_logic_flusher_arbiter (
    .io_inputs_0_valid (TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid     ), //i
    .io_inputs_0_ready (LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready), //o
    .io_output_valid   (LsuPlugin_logic_flusher_arbiter_io_output_valid  ), //o
    .io_output_ready   (LsuPlugin_logic_flusher_arbiter_io_output_ready  ), //i
    .io_chosenOH       (LsuPlugin_logic_flusher_arbiter_io_chosenOH      ), //o
    .clk               (clk                                              ), //i
    .reset             (reset                                            )  //i
  );
  StreamArbiter_3 LsuPlugin_logic_onAddress0_arbiter (
    .io_inputs_0_valid              (LsuPlugin_logic_onAddress0_ls_port_valid                          ), //i
    .io_inputs_0_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_op         (LsuPlugin_logic_onAddress0_ls_port_payload_op[2:0]                ), //i
    .io_inputs_0_payload_address    (LsuPlugin_logic_onAddress0_ls_port_payload_address[31:0]          ), //i
    .io_inputs_0_payload_size       (LsuPlugin_logic_onAddress0_ls_port_payload_size[1:0]              ), //i
    .io_inputs_0_payload_load       (LsuPlugin_logic_onAddress0_ls_port_payload_load                   ), //i
    .io_inputs_0_payload_store      (LsuPlugin_logic_onAddress0_ls_port_payload_store                  ), //i
    .io_inputs_0_payload_atomic     (LsuPlugin_logic_onAddress0_ls_port_payload_atomic                 ), //i
    .io_inputs_0_payload_clean      (LsuPlugin_logic_onAddress0_ls_port_payload_clean                  ), //i
    .io_inputs_0_payload_invalidate (LsuPlugin_logic_onAddress0_ls_port_payload_invalidate             ), //i
    .io_inputs_0_payload_storeId    (LsuPlugin_logic_onAddress0_ls_port_payload_storeId[11:0]          ), //i
    .io_inputs_1_valid              (LsuPlugin_logic_onAddress0_flush_port_valid                       ), //i
    .io_inputs_1_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_op         (LsuPlugin_logic_onAddress0_flush_port_payload_op[2:0]             ), //i
    .io_inputs_1_payload_address    (LsuPlugin_logic_onAddress0_flush_port_payload_address[31:0]       ), //i
    .io_inputs_1_payload_size       (LsuPlugin_logic_onAddress0_flush_port_payload_size[1:0]           ), //i
    .io_inputs_1_payload_load       (LsuPlugin_logic_onAddress0_flush_port_payload_load                ), //i
    .io_inputs_1_payload_store      (LsuPlugin_logic_onAddress0_flush_port_payload_store               ), //i
    .io_inputs_1_payload_atomic     (LsuPlugin_logic_onAddress0_flush_port_payload_atomic              ), //i
    .io_inputs_1_payload_clean      (LsuPlugin_logic_onAddress0_flush_port_payload_clean               ), //i
    .io_inputs_1_payload_invalidate (LsuPlugin_logic_onAddress0_flush_port_payload_invalidate          ), //i
    .io_inputs_1_payload_storeId    (LsuPlugin_logic_onAddress0_flush_port_payload_storeId[11:0]       ), //i
    .io_inputs_2_valid              (LsuPlugin_logic_onAddress0_sb_port_valid                          ), //i
    .io_inputs_2_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready              ), //o
    .io_inputs_2_payload_op         (LsuPlugin_logic_onAddress0_sb_port_payload_op[2:0]                ), //i
    .io_inputs_2_payload_address    (LsuPlugin_logic_onAddress0_sb_port_payload_address[31:0]          ), //i
    .io_inputs_2_payload_size       (LsuPlugin_logic_onAddress0_sb_port_payload_size[1:0]              ), //i
    .io_inputs_2_payload_load       (LsuPlugin_logic_onAddress0_sb_port_payload_load                   ), //i
    .io_inputs_2_payload_store      (LsuPlugin_logic_onAddress0_sb_port_payload_store                  ), //i
    .io_inputs_2_payload_atomic     (LsuPlugin_logic_onAddress0_sb_port_payload_atomic                 ), //i
    .io_inputs_2_payload_clean      (LsuPlugin_logic_onAddress0_sb_port_payload_clean                  ), //i
    .io_inputs_2_payload_invalidate (LsuPlugin_logic_onAddress0_sb_port_payload_invalidate             ), //i
    .io_inputs_2_payload_storeId    (LsuPlugin_logic_onAddress0_sb_port_payload_storeId[11:0]          ), //i
    .io_inputs_3_valid              (LsuPlugin_logic_onAddress0_fromHp_port_valid                      ), //i
    .io_inputs_3_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_3_ready              ), //o
    .io_inputs_3_payload_op         (LsuPlugin_logic_onAddress0_fromHp_port_payload_op[2:0]            ), //i
    .io_inputs_3_payload_address    (LsuPlugin_logic_onAddress0_fromHp_port_payload_address[31:0]      ), //i
    .io_inputs_3_payload_size       (LsuPlugin_logic_onAddress0_fromHp_port_payload_size[1:0]          ), //i
    .io_inputs_3_payload_load       (LsuPlugin_logic_onAddress0_fromHp_port_payload_load               ), //i
    .io_inputs_3_payload_store      (LsuPlugin_logic_onAddress0_fromHp_port_payload_store              ), //i
    .io_inputs_3_payload_atomic     (LsuPlugin_logic_onAddress0_fromHp_port_payload_atomic             ), //i
    .io_inputs_3_payload_clean      (LsuPlugin_logic_onAddress0_fromHp_port_payload_clean              ), //i
    .io_inputs_3_payload_invalidate (LsuPlugin_logic_onAddress0_fromHp_port_payload_invalidate         ), //i
    .io_inputs_3_payload_storeId    (LsuPlugin_logic_onAddress0_fromHp_port_payload_storeId[11:0]      ), //i
    .io_output_valid                (LsuPlugin_logic_onAddress0_arbiter_io_output_valid                ), //o
    .io_output_ready                (LsuPlugin_logic_onAddress0_arbiter_io_output_ready                ), //i
    .io_output_payload_op           (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op[2:0]      ), //o
    .io_output_payload_address      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[31:0]), //o
    .io_output_payload_size         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size[1:0]    ), //o
    .io_output_payload_load         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load         ), //o
    .io_output_payload_store        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store        ), //o
    .io_output_payload_atomic       (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic       ), //o
    .io_output_payload_clean        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean        ), //o
    .io_output_payload_invalidate   (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate   ), //o
    .io_output_payload_storeId      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId[11:0]), //o
    .io_chosen                      (LsuPlugin_logic_onAddress0_arbiter_io_chosen[1:0]                 ), //o
    .io_chosenOH                    (LsuPlugin_logic_onAddress0_arbiter_io_chosenOH[3:0]               ), //o
    .clk                            (clk                                                               ), //i
    .reset                          (reset                                                             )  //i
  );
  StreamArbiter_4 streamArbiter_5 (
    .io_inputs_0_valid                                     (LearnPlugin_logic_buffered_0_valid                                         ), //i
    .io_inputs_0_ready                                     (streamArbiter_5_io_inputs_0_ready                                          ), //o
    .io_inputs_0_payload_pcOnLastSlice                     (LearnPlugin_logic_buffered_0_payload_pcOnLastSlice[31:0]                   ), //i
    .io_inputs_0_payload_pcTarget                          (LearnPlugin_logic_buffered_0_payload_pcTarget[31:0]                        ), //i
    .io_inputs_0_payload_taken                             (LearnPlugin_logic_buffered_0_payload_taken                                 ), //i
    .io_inputs_0_payload_isBranch                          (LearnPlugin_logic_buffered_0_payload_isBranch                              ), //i
    .io_inputs_0_payload_isPush                            (LearnPlugin_logic_buffered_0_payload_isPush                                ), //i
    .io_inputs_0_payload_isPop                             (LearnPlugin_logic_buffered_0_payload_isPop                                 ), //i
    .io_inputs_0_payload_wasWrong                          (LearnPlugin_logic_buffered_0_payload_wasWrong                              ), //i
    .io_inputs_0_payload_badPredictedTarget                (LearnPlugin_logic_buffered_0_payload_badPredictedTarget                    ), //i
    .io_inputs_0_payload_history                           (LearnPlugin_logic_buffered_0_payload_history[11:0]                         ), //i
    .io_inputs_0_payload_uopId                             (LearnPlugin_logic_buffered_0_payload_uopId[15:0]                           ), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]), //i
    .io_inputs_1_valid                                     (LearnPlugin_logic_buffered_1_valid                                         ), //i
    .io_inputs_1_ready                                     (streamArbiter_5_io_inputs_1_ready                                          ), //o
    .io_inputs_1_payload_pcOnLastSlice                     (LearnPlugin_logic_buffered_1_payload_pcOnLastSlice[31:0]                   ), //i
    .io_inputs_1_payload_pcTarget                          (LearnPlugin_logic_buffered_1_payload_pcTarget[31:0]                        ), //i
    .io_inputs_1_payload_taken                             (LearnPlugin_logic_buffered_1_payload_taken                                 ), //i
    .io_inputs_1_payload_isBranch                          (LearnPlugin_logic_buffered_1_payload_isBranch                              ), //i
    .io_inputs_1_payload_isPush                            (LearnPlugin_logic_buffered_1_payload_isPush                                ), //i
    .io_inputs_1_payload_isPop                             (LearnPlugin_logic_buffered_1_payload_isPop                                 ), //i
    .io_inputs_1_payload_wasWrong                          (LearnPlugin_logic_buffered_1_payload_wasWrong                              ), //i
    .io_inputs_1_payload_badPredictedTarget                (LearnPlugin_logic_buffered_1_payload_badPredictedTarget                    ), //i
    .io_inputs_1_payload_history                           (LearnPlugin_logic_buffered_1_payload_history[11:0]                         ), //i
    .io_inputs_1_payload_uopId                             (LearnPlugin_logic_buffered_1_payload_uopId[15:0]                           ), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 (LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 (LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 (LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]), //i
    .io_output_valid                                       (streamArbiter_5_io_output_valid                                            ), //o
    .io_output_ready                                       (LearnPlugin_logic_arbitrated_ready                                         ), //i
    .io_output_payload_pcOnLastSlice                       (streamArbiter_5_io_output_payload_pcOnLastSlice[31:0]                      ), //o
    .io_output_payload_pcTarget                            (streamArbiter_5_io_output_payload_pcTarget[31:0]                           ), //o
    .io_output_payload_taken                               (streamArbiter_5_io_output_payload_taken                                    ), //o
    .io_output_payload_isBranch                            (streamArbiter_5_io_output_payload_isBranch                                 ), //o
    .io_output_payload_isPush                              (streamArbiter_5_io_output_payload_isPush                                   ), //o
    .io_output_payload_isPop                               (streamArbiter_5_io_output_payload_isPop                                    ), //o
    .io_output_payload_wasWrong                            (streamArbiter_5_io_output_payload_wasWrong                                 ), //o
    .io_output_payload_badPredictedTarget                  (streamArbiter_5_io_output_payload_badPredictedTarget                       ), //o
    .io_output_payload_history                             (streamArbiter_5_io_output_payload_history[11:0]                            ), //o
    .io_output_payload_uopId                               (streamArbiter_5_io_output_payload_uopId[15:0]                              ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]   ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]   ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]   ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3   (streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]   ), //o
    .io_chosen                                             (streamArbiter_5_io_chosen                                                  ), //o
    .io_chosenOH                                           (streamArbiter_5_io_chosenOH[1:0]                                           ), //o
    .clk                                                   (clk                                                                        ), //i
    .reset                                                 (reset                                                                      )  //i
  );
  FpuSqrt FpuSqrtPlugin_logic_sqrt (
    .io_input_valid           (FpuSqrtPlugin_logic_sqrt_io_input_valid                ), //i
    .io_input_ready           (FpuSqrtPlugin_logic_sqrt_io_input_ready                ), //o
    .io_input_payload_a       (FpuSqrtPlugin_logic_sqrt_io_input_payload_a[53:0]      ), //i
    .io_output_valid          (FpuSqrtPlugin_logic_sqrt_io_output_valid               ), //o
    .io_output_ready          (1'b0                                                   ), //i
    .io_output_payload_result (FpuSqrtPlugin_logic_sqrt_io_output_payload_result[52:0]), //o
    .io_output_payload_remain (FpuSqrtPlugin_logic_sqrt_io_output_payload_remain[56:0]), //o
    .io_flush                 (execute_ctrl2_down_isReady                             ), //i
    .clk                      (clk                                                    ), //i
    .reset                    (reset                                                  )  //i
  );
  RegFileMem integer_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid       ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address[4:0]), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data[31:0]  ), //i
    .io_writes_0_uopId   (integer_RegFilePlugin_logic_writeMerges_0_bus_uopId[15:0]        ), //i
    .io_writes_1_valid   (integer_RegFilePlugin_logic_writeMerges_1_bus_valid              ), //i
    .io_writes_1_address (integer_RegFilePlugin_logic_writeMerges_1_bus_address[4:0]       ), //i
    .io_writes_1_data    (integer_RegFilePlugin_logic_writeMerges_1_bus_data[31:0]         ), //i
    .io_writes_1_uopId   (integer_RegFilePlugin_logic_writeMerges_1_bus_uopId[15:0]        ), //i
    .io_reads_0_valid    (execute_lane1_bypasser_integer_RS1_port_valid                    ), //i
    .io_reads_0_address  (execute_lane1_bypasser_integer_RS1_port_address[4:0]             ), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[31:0]   ), //o
    .io_reads_1_valid    (execute_lane0_bypasser_integer_RS1_port_valid                    ), //i
    .io_reads_1_address  (execute_lane0_bypasser_integer_RS1_port_address[4:0]             ), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[31:0]   ), //o
    .io_reads_2_valid    (execute_lane0_bypasser_integer_RS2_port_valid                    ), //i
    .io_reads_2_address  (execute_lane0_bypasser_integer_RS2_port_address[4:0]             ), //i
    .io_reads_2_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data[31:0]   ), //o
    .io_reads_3_valid    (execute_lane1_bypasser_integer_RS2_port_valid                    ), //i
    .io_reads_3_address  (execute_lane1_bypasser_integer_RS2_port_address[4:0]             ), //i
    .io_reads_3_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data[31:0]   ), //o
    .clk                 (clk                                                              ), //i
    .reset               (reset                                                            )  //i
  );
  RegFileMem_1 float_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (float_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid       ), //i
    .io_writes_0_address (float_RegFilePlugin_logic_regfile_fpga_io_writes_0_address[4:0]), //i
    .io_writes_0_data    (float_RegFilePlugin_logic_regfile_fpga_io_writes_0_data[63:0]  ), //i
    .io_writes_0_uopId   (float_RegFilePlugin_logic_writeMerges_0_bus_uopId[15:0]        ), //i
    .io_reads_0_valid    (execute_lane0_bypasser_float_RS1_port_valid                    ), //i
    .io_reads_0_address  (execute_lane0_bypasser_float_RS1_port_address[4:0]             ), //i
    .io_reads_0_data     (float_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[63:0]   ), //o
    .io_reads_1_valid    (execute_lane0_bypasser_float_RS2_port_valid                    ), //i
    .io_reads_1_address  (execute_lane0_bypasser_float_RS2_port_address[4:0]             ), //i
    .io_reads_1_data     (float_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[63:0]   ), //o
    .io_reads_2_valid    (execute_lane0_bypasser_float_RS3_port_valid                    ), //i
    .io_reads_2_address  (execute_lane0_bypasser_float_RS3_port_address[4:0]             ), //i
    .io_reads_2_data     (float_RegFilePlugin_logic_regfile_fpga_io_reads_2_data[63:0]   ), //o
    .clk                 (clk                                                            ), //i
    .reset               (reset                                                          )  //i
  );
  always @(*) begin
    case(LsuL1Plugin_logic_refill_read_arbiter_sel)
      1'b0 : _zz_LsuL1Plugin_logic_refill_read_cmdAddress = LsuL1Plugin_logic_refill_slots_0_address[31 : 6];
      default : _zz_LsuL1Plugin_logic_refill_read_cmdAddress = LsuL1Plugin_logic_refill_slots_1_address[31 : 6];
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_bus_read_rsp_payload_id)
      1'b0 : begin
        _zz_LsuL1Plugin_logic_refill_read_rspAddress = LsuL1Plugin_logic_refill_slots_0_address;
        _zz_LsuL1Plugin_logic_refill_read_dirty = LsuL1Plugin_logic_refill_slots_0_dirty;
        _zz_LsuL1Plugin_logic_refill_read_way = LsuL1Plugin_logic_refill_slots_0_way;
      end
      default : begin
        _zz_LsuL1Plugin_logic_refill_read_rspAddress = LsuL1Plugin_logic_refill_slots_1_address;
        _zz_LsuL1Plugin_logic_refill_read_dirty = LsuL1Plugin_logic_refill_slots_1_dirty;
        _zz_LsuL1Plugin_logic_refill_read_way = LsuL1Plugin_logic_refill_slots_1_way;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_writeback_read_arbiter_sel)
      1'b0 : begin
        _zz_LsuL1Plugin_logic_writeback_read_address = LsuL1Plugin_logic_writeback_slots_0_address;
        _zz_LsuL1Plugin_logic_writeback_read_way = LsuL1Plugin_logic_writeback_slots_0_way;
      end
      default : begin
        _zz_LsuL1Plugin_logic_writeback_read_address = LsuL1Plugin_logic_writeback_slots_1_address;
        _zz_LsuL1Plugin_logic_writeback_read_way = LsuL1Plugin_logic_writeback_slots_1_way;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_0_read_rsp;
      default : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_1_read_rsp;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_writeback_write_arbiter_sel)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = LsuL1Plugin_logic_writeback_slots_0_address;
      default : _zz_LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = LsuL1Plugin_logic_writeback_slots_1_address;
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1)
      2'b00 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[63 : 0];
      2'b01 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[127 : 64];
      2'b10 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[191 : 128];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[255 : 192];
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1)
      2'b00 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[63 : 0];
      2'b01 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[127 : 64];
      2'b10 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[191 : 128];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[255 : 192];
    endcase
  end

  always @(*) begin
    case(_zz_60)
      2'b00 : _zz_59 = 2'b00;
      2'b01 : _zz_59 = 2'b01;
      2'b10 : _zz_59 = 2'b01;
      default : _zz_59 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_62)
      3'b000 : _zz_61 = 2'b00;
      3'b001 : _zz_61 = 2'b01;
      3'b010 : _zz_61 = 2'b01;
      3'b011 : _zz_61 = 2'b10;
      3'b100 : _zz_61 = 2'b01;
      3'b101 : _zz_61 = 2'b10;
      3'b110 : _zz_61 = 2'b10;
      default : _zz_61 = 2'b11;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_needFlushSel)
      1'b0 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      end
      default : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_targetWay)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      default : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
    endcase
  end

  always @(*) begin
    case(FetchL1Plugin_logic_bus_rsp_payload_id)
      1'b0 : begin
        _zz_FetchL1Plugin_logic_refill_onRsp_wayToAllocate = FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
        _zz_FetchL1Plugin_logic_refill_onRsp_address = FetchL1Plugin_logic_refill_slots_0_address;
      end
      default : begin
        _zz_FetchL1Plugin_logic_refill_onRsp_wayToAllocate = FetchL1Plugin_logic_refill_slots_1_wayToAllocate;
        _zz_FetchL1Plugin_logic_refill_onRsp_address = FetchL1Plugin_logic_refill_slots_1_address;
      end
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1)
      2'b00 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[63 : 0];
      2'b01 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[127 : 64];
      2'b10 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[191 : 128];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[255 : 192];
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1)
      2'b00 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[63 : 0];
      2'b01 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[127 : 64];
      2'b10 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[191 : 128];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[255 : 192];
    endcase
  end

  always @(*) begin
    case(_zz_64)
      2'b00 : _zz_63 = 2'b00;
      2'b01 : _zz_63 = 2'b01;
      2'b10 : _zz_63 = 2'b01;
      default : _zz_63 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1)
      2'b00 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_0;
      2'b01 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_1;
      2'b10 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_2;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_3;
    endcase
  end

  always @(*) begin
    case(fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE)
      2'b00 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_0;
      2'b01 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_1;
      2'b10 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_2;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_3;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28)
      2'b00 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
      2'b01 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = (_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 | 32'h40000000);
      2'b10 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b111},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = ({{{{{7'h0,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? 7'h3b : 7'h33)} | ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5] == 2'b00) ? 32'h40000000 : 32'h0));
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30)
      3'b000 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b001 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b100;
      3'b010 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b110;
      3'b011 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b111;
      3'b100 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b101 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b110 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b010;
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b011;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28)
      2'b00 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
      2'b01 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = (_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 | 32'h40000000);
      2'b10 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b111},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},7'h13};
      default : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = ({{{{{7'h0,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},(AlignerPlugin_logic_extractors_1_ctx_instruction[12] ? 7'h3b : 7'h33)} | ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5] == 2'b00) ? 32'h40000000 : 32'h0));
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30)
      3'b000 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b001 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b100;
      3'b010 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b110;
      3'b011 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b111;
      3'b100 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b101 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b110 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b010;
      default : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b011;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_1)
      3'b000 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_0;
      3'b001 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      3'b010 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_2;
      3'b011 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      3'b100 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_4;
      3'b101 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_5;
      3'b110 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_6;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_3)
      2'b00 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      2'b01 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      2'b10 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_5;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_5)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4 = LsuPlugin_logic_onCtrl_loadData_splitted_2;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4 = LsuPlugin_logic_onCtrl_loadData_splitted_6;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_7)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6 = LsuPlugin_logic_onCtrl_loadData_splitted_3;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6 = LsuPlugin_logic_onCtrl_loadData_splitted_7;
    endcase
  end

  always @(*) begin
    case(_zz_67)
      3'b000 : _zz_66 = _zz_49;
      3'b001 : _zz_66 = _zz_50;
      3'b010 : _zz_66 = _zz_51;
      3'b011 : _zz_66 = _zz_52;
      3'b100 : _zz_66 = _zz_53;
      3'b101 : _zz_66 = _zz_54;
      3'b110 : _zz_66 = _zz_55;
      default : _zz_66 = _zz_56;
    endcase
  end

  always @(*) begin
    case(_zz_69)
      3'b000 : _zz_68 = _zz_49;
      3'b001 : _zz_68 = _zz_50;
      3'b010 : _zz_68 = _zz_51;
      3'b011 : _zz_68 = _zz_52;
      3'b100 : _zz_68 = _zz_53;
      3'b101 : _zz_68 = _zz_54;
      3'b110 : _zz_68 = _zz_55;
      default : _zz_68 = _zz_56;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_candidates_1_age_1)
      1'b0 : _zz_DispatchPlugin_logic_candidates_1_age = 1'b0;
      default : _zz_DispatchPlugin_logic_candidates_1_age = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_candidates_2_age_1)
      2'b00 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b00;
      2'b01 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b01;
      2'b10 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b01;
      default : _zz_DispatchPlugin_logic_candidates_2_age = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_slotsFeeds_fit_1)
      2'b00 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b00;
      2'b01 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b01;
      2'b10 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b01;
      default : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b10;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      1'b0 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = TrapPlugin_logic_harts_0_crsPorts_read_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = CsrRamPlugin_csrMapper_read_address;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_candidatesCount_1)
      3'b000 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b00;
      3'b001 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b010 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b011 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      3'b100 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b101 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      3'b110 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      default : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b11;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1)
      2'b00 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b00;
      2'b01 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b01;
      2'b10 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b01;
      default : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl4_down_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl4_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl4_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl4_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_up_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl5_up_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_up_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl5_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl5_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl5_up_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl4_up_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl4_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl4_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl4_up_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl3_up_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl3_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl3_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl3_up_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl2_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl2_up_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl2_up_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_down_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl5_down_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl5_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl5_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl5_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl3_down_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl3_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl3_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl3_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : execute_ctrl2_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : execute_ctrl2_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : execute_ctrl2_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE)
      FpuRoundMode_RNE : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "RMM";
      default : FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuPackerPlugin_logic_pip_node_2_s0_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuPackerPlugin_logic_pip_node_2_s0_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuPackerPlugin_logic_pip_node_2_s0_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE)
      FpuRoundMode_RNE : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "RMM";
      default : FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_1_s0_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuPackerPlugin_logic_pip_node_1_s0_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuPackerPlugin_logic_pip_node_1_s0_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuPackerPlugin_logic_pip_node_1_s0_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE)
      FpuRoundMode_RNE : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RMM";
      default : FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_0_s0_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "RNE";
      FpuRoundMode_RTZ : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "RTZ";
      FpuRoundMode_RDN : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "RDN";
      FpuRoundMode_RUP : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "RUP";
      FpuRoundMode_RMM : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "RMM";
      default : execute_ctrl2_down_FpuUtils_ROUNDING_lane0_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "RMM";
      default : FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "RMM";
      default : FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "RMM";
      default : FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "RMM";
      default : FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RMM";
      default : FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(FpuUnpackerPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuUnpackerPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuUnpackerPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuUnpackerPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuUnpackerPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuUnpackerPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuUnpackerPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuUnpackerPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddPlugin_logic_addPort_cmd_rs1_mode)
      FloatMode_ZERO : FpuAddPlugin_logic_addPort_cmd_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddPlugin_logic_addPort_cmd_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddPlugin_logic_addPort_cmd_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddPlugin_logic_addPort_cmd_rs1_mode_string = "NORMAL";
      default : FpuAddPlugin_logic_addPort_cmd_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddPlugin_logic_addPort_cmd_rs2_mode)
      FloatMode_ZERO : FpuAddPlugin_logic_addPort_cmd_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddPlugin_logic_addPort_cmd_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuAddPlugin_logic_addPort_cmd_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddPlugin_logic_addPort_cmd_rs2_mode_string = "NORMAL";
      default : FpuAddPlugin_logic_addPort_cmd_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddPlugin_logic_addPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddPlugin_logic_addPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddPlugin_logic_addPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddPlugin_logic_addPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddPlugin_logic_addPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "RMM";
      default : FpuAddPlugin_logic_addPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuMulPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuMulPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuMulPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuMulPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuMulPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuMulPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuMulPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuMulPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuMulPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuSqrtPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuSqrtPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuSqrtPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuSqrtPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuSqrtPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuSqrtPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuSqrtPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuSqrtPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuSqrtPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuSqrtPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuSqrtPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuSqrtPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuXxPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuXxPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuXxPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuXxPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuXxPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuXxPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuXxPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuXxPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuXxPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuXxPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuXxPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuXxPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuDivPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuDivPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuDivPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuDivPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuDivPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuDivPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuDivPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuDivPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuDivPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuDivPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuDivPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuDivPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_addPort_cmd_rs1_mode)
      FloatMode_ZERO : FpuMulPlugin_logic_addPort_cmd_rs1_mode_string = "ZERO  ";
      FloatMode_INF : FpuMulPlugin_logic_addPort_cmd_rs1_mode_string = "INF   ";
      FloatMode_NAN : FpuMulPlugin_logic_addPort_cmd_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuMulPlugin_logic_addPort_cmd_rs1_mode_string = "NORMAL";
      default : FpuMulPlugin_logic_addPort_cmd_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_addPort_cmd_rs2_mode)
      FloatMode_ZERO : FpuMulPlugin_logic_addPort_cmd_rs2_mode_string = "ZERO  ";
      FloatMode_INF : FpuMulPlugin_logic_addPort_cmd_rs2_mode_string = "INF   ";
      FloatMode_NAN : FpuMulPlugin_logic_addPort_cmd_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuMulPlugin_logic_addPort_cmd_rs2_mode_string = "NORMAL";
      default : FpuMulPlugin_logic_addPort_cmd_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_addPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuMulPlugin_logic_addPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuMulPlugin_logic_addPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuMulPlugin_logic_addPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_addPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "RMM";
      default : FpuMulPlugin_logic_addPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_packPort_cmd_value_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_packPort_cmd_value_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : FpuAddSharedPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuAddSharedPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : FpuAddSharedPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_packPort_cmd_roundMode)
      FpuRoundMode_RNE : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "RMM";
      default : FpuAddSharedPlugin_logic_packPort_cmd_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode)
      FloatMode_ZERO : FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string = "ZERO  ";
      FloatMode_INF : FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string = "INF   ";
      FloatMode_NAN : FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string = "NORMAL";
      default : FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode)
      FloatMode_ZERO : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "ZERO  ";
      FloatMode_INF : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "INF   ";
      FloatMode_NAN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "NORMAL";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1)
      FloatMode_ZERO : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string = "NORMAL";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode)
      FloatMode_ZERO : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "ZERO  ";
      FloatMode_INF : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "INF   ";
      FloatMode_NAN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "NORMAL";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1)
      FloatMode_ZERO : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string = "NORMAL";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE)
      FpuRoundMode_RNE : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "RMM";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1)
      FpuRoundMode_RNE : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "RMM";
      default : _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1)
      FpuRoundMode_RNE : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "RNE";
      FpuRoundMode_RTZ : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "RTZ";
      FpuRoundMode_RDN : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "RDN";
      FpuRoundMode_RUP : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "RUP";
      FpuRoundMode_RMM : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "RMM";
      default : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1_string = "???";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_ls_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_flush_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_sb_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_sb_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_fromHp_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_fromHp_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_0_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_0_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_0_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_0_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_0_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_1_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_1_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_1_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_1_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_1_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_1_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_2_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_2_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_2_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_2_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_2_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_2_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_3_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_3_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_3_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_3_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_3_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_3_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_4_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_4_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_4_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_4_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_4_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_4_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPackerPlugin_logic_s0_remapped_5_mode)
      FloatMode_ZERO : FpuPackerPlugin_logic_s0_remapped_5_mode_string = "ZERO  ";
      FloatMode_INF : FpuPackerPlugin_logic_s0_remapped_5_mode_string = "INF   ";
      FloatMode_NAN : FpuPackerPlugin_logic_s0_remapped_5_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuPackerPlugin_logic_s0_remapped_5_mode_string = "NORMAL";
      default : FpuPackerPlugin_logic_s0_remapped_5_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode)
      FloatMode_ZERO : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "ZERO  ";
      FloatMode_INF : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "INF   ";
      FloatMode_NAN : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "NORMAL";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1)
      FloatMode_ZERO : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string = "NORMAL";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE)
      FpuRoundMode_RNE : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "RMM";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1)
      FpuRoundMode_RNE : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "RMM";
      default : _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2)
      FloatMode_ZERO : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string = "ZERO  ";
      FloatMode_INF : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string = "INF   ";
      FloatMode_NAN : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string = "NAN   ";
      FloatMode_NORMAL : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string = "NORMAL";
      default : _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuMulPlugin_logic_onPack_mode)
      FloatMode_ZERO : FpuMulPlugin_logic_onPack_mode_string = "ZERO  ";
      FloatMode_INF : FpuMulPlugin_logic_onPack_mode_string = "INF   ";
      FloatMode_NAN : FpuMulPlugin_logic_onPack_mode_string = "NAN   ";
      FloatMode_NORMAL : FpuMulPlugin_logic_onPack_mode_string = "NORMAL";
      default : FpuMulPlugin_logic_onPack_mode_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuXxPlugin_logic_packPort_cmd_format)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_FpuXxPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_FpuXxPlugin_logic_packPort_cmd_format_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_FpuXxPlugin_logic_packPort_cmd_format_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2)
      FpuFormat_FpuCmpPlugin_logic_f32_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2_string = "FpuCmpPlugin_logic_f32_1";
      FpuFormat_FpuCmpPlugin_logic_f64_1 : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2_string = "FpuCmpPlugin_logic_f64_1";
      default : _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0)
      FpuCmpFloatOp_MIN_MAX : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "SGNJ   ";
      default : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1)
      FpuCmpFloatOp_MIN_MAX : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1_string = "SGNJ   ";
      default : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2)
      FpuCmpFloatOp_MIN_MAX : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2_string = "MIN_MAX";
      FpuCmpFloatOp_SGNJ : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2_string = "SGNJ   ";
      default : _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "ZERO ";
      default : _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "?????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateReg_string = "IDLE      ";
      LsuPlugin_logic_flusher_SB_DRAIN : LsuPlugin_logic_flusher_stateReg_string = "SB_DRAIN  ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateReg_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateReg_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateNext)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateNext_string = "IDLE      ";
      LsuPlugin_logic_flusher_SB_DRAIN : LsuPlugin_logic_flusher_stateNext_string = "SB_DRAIN  ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateNext_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateNext_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "COMPUTE    ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateNext)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "COMPUTE    ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "???????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateReg_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateReg_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateNext)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateNext_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateNext_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    BtbPlugin_logic_ras_ptr_pop_aheadValue = BtbPlugin_logic_ras_ptr_pop;
    BtbPlugin_logic_ras_ptr_pop_aheadValue = (_zz_BtbPlugin_logic_ras_ptr_pop_aheadValue - _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3);
  end

  assign execute_ctrl4_down_RD_ENABLE_lane1 = execute_ctrl4_RD_ENABLE_lane1_bypass;
  always @(*) begin
    execute_ctrl4_RD_ENABLE_lane1_bypass = execute_ctrl4_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l306_9) begin
      execute_ctrl4_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_LANE_SEL_lane1 = execute_ctrl4_LANE_SEL_lane1_bypass;
  always @(*) begin
    execute_ctrl4_LANE_SEL_lane1_bypass = execute_ctrl4_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l306_9) begin
      execute_ctrl4_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_RD_ENABLE_lane1 = execute_ctrl3_RD_ENABLE_lane1_bypass;
  always @(*) begin
    execute_ctrl3_RD_ENABLE_lane1_bypass = execute_ctrl3_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l306_8) begin
      execute_ctrl3_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LANE_SEL_lane1 = execute_ctrl3_LANE_SEL_lane1_bypass;
  always @(*) begin
    execute_ctrl3_LANE_SEL_lane1_bypass = execute_ctrl3_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l306_8) begin
      execute_ctrl3_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_RD_ENABLE_lane1 = execute_ctrl2_RD_ENABLE_lane1_bypass;
  always @(*) begin
    execute_ctrl2_RD_ENABLE_lane1_bypass = execute_ctrl2_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l306_7) begin
      execute_ctrl2_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_LANE_SEL_lane1 = execute_ctrl2_LANE_SEL_lane1_bypass;
  always @(*) begin
    execute_ctrl2_LANE_SEL_lane1_bypass = execute_ctrl2_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l306_7) begin
      execute_ctrl2_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_RD_ENABLE_lane1 = execute_ctrl1_RD_ENABLE_lane1_bypass;
  always @(*) begin
    execute_ctrl1_RD_ENABLE_lane1_bypass = execute_ctrl1_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l306_6) begin
      execute_ctrl1_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_LANE_SEL_lane1 = execute_ctrl1_LANE_SEL_lane1_bypass;
  always @(*) begin
    execute_ctrl1_LANE_SEL_lane1_bypass = execute_ctrl1_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l306_6) begin
      execute_ctrl1_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_RD_ENABLE_lane1 = execute_ctrl0_RD_ENABLE_lane1_bypass;
  always @(*) begin
    execute_ctrl0_RD_ENABLE_lane1_bypass = execute_ctrl0_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l306_5) begin
      execute_ctrl0_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_LANE_SEL_lane1 = execute_ctrl0_LANE_SEL_lane1_bypass;
  always @(*) begin
    execute_ctrl0_LANE_SEL_lane1_bypass = execute_ctrl0_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l306_5) begin
      execute_ctrl0_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_integer_RS2_lane1 = execute_ctrl3_integer_RS2_lane1_bypass;
  assign execute_ctrl2_down_integer_RS2_lane1 = execute_ctrl2_integer_RS2_lane1_bypass;
  assign execute_ctrl3_down_integer_RS1_lane1 = execute_ctrl3_integer_RS1_lane1_bypass;
  assign execute_ctrl2_down_integer_RS1_lane1 = execute_ctrl2_integer_RS1_lane1_bypass;
  assign execute_ctrl4_down_RD_ENABLE_lane0 = execute_ctrl4_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl4_RD_ENABLE_lane0_bypass = execute_ctrl4_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_LANE_SEL_lane0 = execute_ctrl4_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LANE_SEL_lane0_bypass = execute_ctrl4_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_RD_ENABLE_lane0 = execute_ctrl3_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl3_RD_ENABLE_lane0_bypass = execute_ctrl3_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LANE_SEL_lane0 = execute_ctrl3_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LANE_SEL_lane0_bypass = execute_ctrl3_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_RD_ENABLE_lane0 = execute_ctrl2_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl2_RD_ENABLE_lane0_bypass = execute_ctrl2_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_LANE_SEL_lane0 = execute_ctrl2_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl2_LANE_SEL_lane0_bypass = execute_ctrl2_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_RD_ENABLE_lane0 = execute_ctrl1_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl1_RD_ENABLE_lane0_bypass = execute_ctrl1_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_LANE_SEL_lane0 = execute_ctrl1_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl1_LANE_SEL_lane0_bypass = execute_ctrl1_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_RD_ENABLE_lane0 = execute_ctrl0_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl0_RD_ENABLE_lane0_bypass = execute_ctrl0_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_LANE_SEL_lane0 = execute_ctrl0_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl0_LANE_SEL_lane0_bypass = execute_ctrl0_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_integer_RS2_lane0 = execute_ctrl3_integer_RS2_lane0_bypass;
  assign execute_ctrl2_down_integer_RS2_lane0 = execute_ctrl2_integer_RS2_lane0_bypass;
  assign execute_ctrl3_down_integer_RS1_lane0 = execute_ctrl3_integer_RS1_lane0_bypass;
  assign execute_ctrl2_down_integer_RS1_lane0 = execute_ctrl2_integer_RS1_lane0_bypass;
  always @(*) begin
    _zz_1 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_fault;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_fault_1 = _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1[0];
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_target;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_target_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_pc : 32'h0);
    end
  end

  assign decode_ctrls_1_down_LANE_SEL_1 = decode_ctrls_1_LANE_SEL_1_bypass;
  always @(*) begin
    decode_ctrls_1_LANE_SEL_1_bypass = decode_ctrls_1_up_LANE_SEL_1;
    if(decode_logic_flushes_1_onLanes_1_doIt) begin
      decode_ctrls_1_LANE_SEL_1_bypass = 1'b0;
    end
  end

  assign decode_ctrls_1_down_LANE_SEL_0 = decode_ctrls_1_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_1_LANE_SEL_0_bypass = decode_ctrls_1_up_LANE_SEL_0;
    if(decode_logic_flushes_1_onLanes_0_doIt) begin
      decode_ctrls_1_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign decode_ctrls_0_down_LANE_SEL_1 = decode_ctrls_0_LANE_SEL_1_bypass;
  always @(*) begin
    decode_ctrls_0_LANE_SEL_1_bypass = decode_ctrls_0_up_LANE_SEL_1;
    if(decode_logic_flushes_0_onLanes_1_doIt) begin
      decode_ctrls_0_LANE_SEL_1_bypass = 1'b0;
    end
  end

  assign decode_ctrls_0_down_LANE_SEL_0 = decode_ctrls_0_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_0_LANE_SEL_0_bypass = decode_ctrls_0_up_LANE_SEL_0;
    if(decode_logic_flushes_0_onLanes_0_doIt) begin
      decode_ctrls_0_LANE_SEL_0_bypass = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[5] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6_1 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5);
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[4] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4);
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[3] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3);
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[2] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2);
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[1] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1);
  end

  always @(*) begin
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
    execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[0] ? _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 : execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0);
  end

  always @(*) begin
    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 = _zz_when_Utils_l1585;
    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 = (_zz_when_Utils_l1585_17[3] ? _zz__zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 : _zz_when_Utils_l1585);
  end

  always @(*) begin
    _zz_when_Utils_l1585 = _zz_when_Utils_l1585_1;
    _zz_when_Utils_l1585 = (_zz_when_Utils_l1585_17[2] ? _zz__zz_when_Utils_l1585 : _zz_when_Utils_l1585_1);
  end

  always @(*) begin
    _zz_when_Utils_l1585_1 = _zz_when_Utils_l1585_2;
    _zz_when_Utils_l1585_1 = (_zz_when_Utils_l1585_17[1] ? _zz__zz_when_Utils_l1585_1 : _zz_when_Utils_l1585_2);
  end

  always @(*) begin
    _zz_when_Utils_l1585_2 = _zz_when_Utils_l1585_16;
    _zz_when_Utils_l1585_2 = (_zz_when_Utils_l1585_17[0] ? _zz__zz_when_Utils_l1585_2 : _zz_when_Utils_l1585_16);
  end

  assign execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl11_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl8_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl7_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl5_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl4_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl3_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl3_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  assign execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign decode_ctrls_1_down_TRAP_1 = decode_ctrls_1_TRAP_1_bypass;
  always @(*) begin
    decode_ctrls_1_TRAP_1_bypass = decode_ctrls_1_up_TRAP_1;
    if(when_DecoderPlugin_l229_1) begin
      decode_ctrls_1_TRAP_1_bypass = 1'b1;
    end
  end

  assign decode_ctrls_1_down_TRAP_0 = decode_ctrls_1_TRAP_0_bypass;
  always @(*) begin
    decode_ctrls_1_TRAP_0_bypass = decode_ctrls_1_up_TRAP_0;
    if(when_DecoderPlugin_l229) begin
      decode_ctrls_1_TRAP_0_bypass = 1'b1;
    end
  end

  assign execute_ctrl2_down_COMPLETED_lane0 = execute_ctrl2_COMPLETED_lane0_bypass;
  assign execute_ctrl8_down_COMPLETED_lane0 = execute_ctrl8_COMPLETED_lane0_bypass;
  assign execute_ctrl5_down_COMPLETED_lane0 = execute_ctrl5_COMPLETED_lane0_bypass;
  assign execute_ctrl3_down_COMPLETED_lane0 = execute_ctrl3_COMPLETED_lane0_bypass;
  assign execute_ctrl11_down_COMPLETED_lane0 = execute_ctrl11_COMPLETED_lane0_bypass;
  assign execute_ctrl7_down_COMPLETED_lane0 = execute_ctrl7_COMPLETED_lane0_bypass;
  assign execute_ctrl4_down_COMPLETED_lane0 = execute_ctrl4_COMPLETED_lane0_bypass;
  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_shifter_4 = late1_BranchPlugin_logic_jumpLogic_history_shifter_3;
    if(when_BranchPlugin_l218_3) begin
      late1_BranchPlugin_logic_jumpLogic_history_shifter_4 = _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_shifter_3 = late1_BranchPlugin_logic_jumpLogic_history_shifter_2;
    if(when_BranchPlugin_l213_11) begin
      late1_BranchPlugin_logic_jumpLogic_history_shifter_3 = _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_shifter_2 = late1_BranchPlugin_logic_jumpLogic_history_shifter_1;
    if(when_BranchPlugin_l213_10) begin
      late1_BranchPlugin_logic_jumpLogic_history_shifter_2 = _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_shifter_1 = late1_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l213_9) begin
      late1_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_late1_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_shifter_4 = late0_BranchPlugin_logic_jumpLogic_history_shifter_3;
    if(when_BranchPlugin_l218_2) begin
      late0_BranchPlugin_logic_jumpLogic_history_shifter_4 = _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_shifter_3 = late0_BranchPlugin_logic_jumpLogic_history_shifter_2;
    if(when_BranchPlugin_l213_8) begin
      late0_BranchPlugin_logic_jumpLogic_history_shifter_3 = _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_shifter_2 = late0_BranchPlugin_logic_jumpLogic_history_shifter_1;
    if(when_BranchPlugin_l213_7) begin
      late0_BranchPlugin_logic_jumpLogic_history_shifter_2 = _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_shifter_1 = late0_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l213_6) begin
      late0_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_late0_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  assign execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX = execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX;
  assign execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF = execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_UF;
  assign execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF = execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_OF;
  assign execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ = execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_DZ;
  assign execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV = execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NV;
  assign execute_ctrl4_down_COMPLETED_lane1 = execute_ctrl4_COMPLETED_lane1_bypass;
  assign execute_ctrl2_down_COMPLETED_lane1 = execute_ctrl2_COMPLETED_lane1_bypass;
  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_shifter_4 = early1_BranchPlugin_logic_jumpLogic_history_shifter_3;
    if(when_BranchPlugin_l218_1) begin
      early1_BranchPlugin_logic_jumpLogic_history_shifter_4 = _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_shifter_3 = early1_BranchPlugin_logic_jumpLogic_history_shifter_2;
    if(when_BranchPlugin_l213_5) begin
      early1_BranchPlugin_logic_jumpLogic_history_shifter_3 = _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_shifter_2 = early1_BranchPlugin_logic_jumpLogic_history_shifter_1;
    if(when_BranchPlugin_l213_4) begin
      early1_BranchPlugin_logic_jumpLogic_history_shifter_2 = _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_shifter_1 = early1_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l213_3) begin
      early1_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_early1_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_4 = early0_BranchPlugin_logic_jumpLogic_history_shifter_3;
    if(when_BranchPlugin_l218) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_4 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_3 = early0_BranchPlugin_logic_jumpLogic_history_shifter_2;
    if(when_BranchPlugin_l213_2) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_3 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
    if(when_BranchPlugin_l213_1) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_2 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = early0_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l213) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter = _zz_when_Utils_l1585_3;
    _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter = (FpuPackerPlugin_logic_s1_subnormal_manShift[5] ? _zz__zz_FpuPackerPlugin_logic_s1_subnormal_manShifter : _zz_when_Utils_l1585_3);
  end

  always @(*) begin
    _zz_when_Utils_l1585_3 = _zz_when_Utils_l1585_4;
    _zz_when_Utils_l1585_3 = (FpuPackerPlugin_logic_s1_subnormal_manShift[4] ? _zz__zz_when_Utils_l1585_3 : _zz_when_Utils_l1585_4);
  end

  always @(*) begin
    _zz_when_Utils_l1585_4 = _zz_when_Utils_l1585_5;
    _zz_when_Utils_l1585_4 = (FpuPackerPlugin_logic_s1_subnormal_manShift[3] ? _zz__zz_when_Utils_l1585_4 : _zz_when_Utils_l1585_5);
  end

  always @(*) begin
    _zz_when_Utils_l1585_5 = _zz_when_Utils_l1585_6;
    _zz_when_Utils_l1585_5 = (FpuPackerPlugin_logic_s1_subnormal_manShift[2] ? _zz__zz_when_Utils_l1585_5 : _zz_when_Utils_l1585_6);
  end

  always @(*) begin
    _zz_when_Utils_l1585_6 = _zz_when_Utils_l1585_7;
    _zz_when_Utils_l1585_6 = (FpuPackerPlugin_logic_s1_subnormal_manShift[1] ? _zz__zz_when_Utils_l1585_6 : _zz_when_Utils_l1585_7);
  end

  always @(*) begin
    _zz_when_Utils_l1585_7 = _zz_when_Utils_l1585_15;
    _zz_when_Utils_l1585_7 = (FpuPackerPlugin_logic_s1_subnormal_manShift[0] ? _zz__zz_when_Utils_l1585_7 : _zz_when_Utils_l1585_15);
  end

  assign execute_ctrl4_down_COMMIT_lane0 = execute_ctrl4_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl4_COMMIT_lane0_bypass = execute_ctrl4_up_COMMIT_lane0;
    if(when_LsuPlugin_l865) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_COMMIT_lane0_bypass = 1'b0;
      end
    end
  end

  assign execute_ctrl4_down_TRAP_lane0 = execute_ctrl4_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl4_TRAP_lane0_bypass = execute_ctrl4_up_TRAP_lane0;
    if(when_LsuPlugin_l865) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_TRAP_lane0_bypass = 1'b1;
      end
    end
  end

  assign execute_ctrl4_down_LsuL1_SEL_lane0 = execute_ctrl4_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LsuL1_SEL_lane0_bypass = execute_ctrl4_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l546_1) begin
      execute_ctrl4_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LsuL1_SEL_lane0 = execute_ctrl3_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LsuL1_SEL_lane0_bypass = execute_ctrl3_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l546) begin
      execute_ctrl3_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(LsuPlugin_logic_storeBuffer_push_valid) begin
      _zz_2 = 1'b1;
    end
  end

  assign execute_ctrl2_down_COMMIT_lane0 = execute_ctrl2_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl2_COMMIT_lane0_bypass = execute_ctrl2_up_COMMIT_lane0;
    if(when_EnvPlugin_l119) begin
      if(when_EnvPlugin_l123) begin
        execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
      end
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
            end
          end
        end
      end
    endcase
  end

  assign execute_ctrl2_down_TRAP_lane0 = execute_ctrl2_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl2_TRAP_lane0_bypass = execute_ctrl2_up_TRAP_lane0;
    if(when_EnvPlugin_l119) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_TRAP_lane0_bypass = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                execute_ctrl2_TRAP_lane0_bypass = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter = _zz_when_Utils_l1585_8;
    _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[6] ? _zz__zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter : _zz_when_Utils_l1585_8);
  end

  always @(*) begin
    _zz_when_Utils_l1585_8 = _zz_when_Utils_l1585_9;
    _zz_when_Utils_l1585_8 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[5] ? _zz__zz_when_Utils_l1585_8 : _zz_when_Utils_l1585_9);
  end

  always @(*) begin
    _zz_when_Utils_l1585_9 = _zz_when_Utils_l1585_10;
    _zz_when_Utils_l1585_9 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[4] ? _zz__zz_when_Utils_l1585_9 : _zz_when_Utils_l1585_10);
  end

  always @(*) begin
    _zz_when_Utils_l1585_10 = _zz_when_Utils_l1585_11;
    _zz_when_Utils_l1585_10 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[3] ? _zz__zz_when_Utils_l1585_10 : _zz_when_Utils_l1585_11);
  end

  always @(*) begin
    _zz_when_Utils_l1585_11 = _zz_when_Utils_l1585_12;
    _zz_when_Utils_l1585_11 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[2] ? _zz__zz_when_Utils_l1585_11 : _zz_when_Utils_l1585_12);
  end

  always @(*) begin
    _zz_when_Utils_l1585_12 = _zz_when_Utils_l1585_13;
    _zz_when_Utils_l1585_12 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[1] ? _zz__zz_when_Utils_l1585_12 : _zz_when_Utils_l1585_13);
  end

  always @(*) begin
    _zz_when_Utils_l1585_13 = _zz_when_Utils_l1585_14;
    _zz_when_Utils_l1585_13 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[0] ? _zz__zz_when_Utils_l1585_13 : _zz_when_Utils_l1585_14);
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(BtbPlugin_logic_ras_write_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(GSharePlugin_logic_mem_writes_0_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(FetchL1Plugin_logic_plru_write_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(FetchL1Plugin_logic_banks_1_write_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(FetchL1Plugin_logic_banks_0_write_valid) begin
      _zz_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_8 = 1'b0;
    if(PrefetcherRptPlugin_logic_storage_write_valid) begin
      _zz_8 = 1'b1;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  always @(*) begin
    _zz_9 = 1'b0;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      _zz_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_10 = 1'b0;
    if(LsuL1Plugin_logic_shared_write_valid) begin
      _zz_10 = 1'b1;
    end
  end

  assign AlignerPlugin_api_singleFetch = 1'b0;
  assign AlignerPlugin_api_haltIt = 1'b0;
  always @(*) begin
    DispatchPlugin_api_haltDispatch = 1'b0;
    if(_zz_25) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
    if(LsuPlugin_logic_storeBuffer_holdHart_waitIt) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
  end

  assign CsrRamPlugin_api_holdRead = 1'b0;
  assign CsrRamPlugin_api_holdWrite = 1'b0;
  assign PrivilegedPlugin_api_harts_0_allowInterrupts = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowEbreakException = 1'b1;
  always @(*) begin
    PrivilegedPlugin_api_harts_0_fpuEnable = 1'b0;
    if(when_PrivilegedPlugin_l549) begin
      PrivilegedPlugin_api_harts_0_fpuEnable = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_redo = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
              TrapPlugin_api_harts_0_redo = 1'b1;
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_api_harts_0_askWake = 1'b0;
    if(when_TrapPlugin_l226) begin
      TrapPlugin_api_harts_0_askWake = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_rvTrap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_api_harts_0_rvTrap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuCsrPlugin_api_gotDirty = 1'b0;
    if(when_FpuCsrPlugin_l61) begin
      FpuCsrPlugin_api_gotDirty = 1'b1;
    end
    if(when_CsrAccessPlugin_l346_7) begin
      FpuCsrPlugin_api_gotDirty = 1'b1;
    end
  end

  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 & execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 | execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 ^ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        early0_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign early0_IntAluPlugin_logic_alu_result = (_zz_early0_IntAluPlugin_logic_alu_result | _zz_early0_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0 = early0_IntAluPlugin_logic_alu_result;
  assign early0_IntAluPlugin_logic_wb_valid = execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  assign early0_IntAluPlugin_logic_wb_payload = execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  assign early0_BarrelShifterPlugin_logic_shift_amplitude = _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  assign early0_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0);
  assign early0_BarrelShifterPlugin_logic_shift_shifted = _zz_early0_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign early0_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_patched : early0_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = early0_BarrelShifterPlugin_logic_shift_patched;
  assign early0_BarrelShifterPlugin_logic_wb_valid = execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  assign early0_BarrelShifterPlugin_logic_wb_payload = execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  always @(*) begin
    LsuL1_ackUnlock = 1'b0;
    if(LsuPlugin_logic_onCtrl_io_cmdSent) begin
      LsuL1_ackUnlock = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_address = 7'bxxxxxxx;
    LsuL1Plugin_logic_banksWrite_address = {LsuL1Plugin_logic_refill_read_rspAddress[11 : 6],LsuL1Plugin_logic_refill_read_wordIndex};
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 5];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeData = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeData = LsuL1Plugin_logic_bus_read_rsp_payload_data;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeData[63 : 0] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
      LsuL1Plugin_logic_banksWrite_writeData[127 : 64] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
      LsuL1Plugin_logic_banksWrite_writeData[191 : 128] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
      LsuL1Plugin_logic_banksWrite_writeData[255 : 192] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeMask = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeMask = 32'hffffffff;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeMask = 32'h0;
      if(_zz_24[0]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[7 : 0] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
      if(_zz_24[1]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[15 : 8] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
      if(_zz_24[2]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[23 : 16] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
      if(_zz_24[3]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[31 : 24] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
        LsuL1Plugin_logic_banksWrite_writeMask = 32'h0;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_mask = 2'b00;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_mask[LsuL1Plugin_logic_refill_read_way] = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_mask = LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) begin
        LsuL1Plugin_logic_waysWrite_mask = 2'b00;
      end
    end
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_waysWrite_mask = 2'b11;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_refill_read_rspAddress[11 : 6];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    end
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_address = LsuL1Plugin_logic_refill_read_rspAddress[31 : 12];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_address = _zz_LsuL1Plugin_logic_waysWrite_tag_address;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_fault = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_fault = LsuL1Plugin_logic_refill_read_faulty;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_fault = _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
    end
  end

  assign LsuL1Plugin_logic_waysWrite_valid = (|LsuL1Plugin_logic_waysWrite_mask);
  assign LsuL1Plugin_logic_banks_0_write_valid = LsuL1Plugin_logic_banksWrite_mask[0];
  assign LsuL1Plugin_logic_banks_0_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_0_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_0_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_0_read_rsp = LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_banks_1_write_valid = LsuL1Plugin_logic_banksWrite_mask[1];
  assign LsuL1Plugin_logic_banks_1_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_1_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_1_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_1_read_rsp = LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  assign _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = LsuL1Plugin_logic_shared_mem_spinal_port1;
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1[0 : 0];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_dirty = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[2 : 1];
  always @(*) begin
    LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        case(LsuL1Plugin_logic_bus_read_rsp_payload_id)
          1'b0 : begin
            LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
  end

  assign LsuL1Plugin_logic_refill_slots_0_loadedDone = (LsuL1Plugin_logic_refill_slots_0_loadedCounter == 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_free = ((! LsuL1Plugin_logic_refill_slots_0_valid) && 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_fire = ((! execute_freeze_valid) && LsuL1Plugin_logic_refill_slots_0_loadedDone);
  always @(*) begin
    LsuL1Plugin_logic_refill_slots_1_loadedSet = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        case(LsuL1Plugin_logic_bus_read_rsp_payload_id)
          1'b0 : begin
          end
          default : begin
            LsuL1Plugin_logic_refill_slots_1_loadedSet = 1'b1;
          end
        endcase
      end
    end
  end

  assign LsuL1Plugin_logic_refill_slots_1_loadedDone = (LsuL1Plugin_logic_refill_slots_1_loadedCounter == 1'b1);
  assign LsuL1Plugin_logic_refill_slots_1_free = ((! LsuL1Plugin_logic_refill_slots_1_valid) && 1'b1);
  assign LsuL1Plugin_logic_refill_slots_1_fire = ((! execute_freeze_valid) && LsuL1Plugin_logic_refill_slots_1_loadedDone);
  assign _zz_LsuL1Plugin_logic_refill_free = {LsuL1Plugin_logic_refill_slots_1_free,LsuL1Plugin_logic_refill_slots_0_free};
  assign LsuL1Plugin_logic_refill_free = {_zz_LsuL1Plugin_logic_refill_free_1[1],LsuL1Plugin_logic_refill_slots_0_free};
  assign LsuL1Plugin_logic_refill_full = (&{(! LsuL1Plugin_logic_refill_slots_1_free),(! LsuL1Plugin_logic_refill_slots_0_free)});
  assign when_LsuL1Plugin_l377 = (LsuL1Plugin_logic_refill_push_valid && LsuL1Plugin_logic_refill_free[0]);
  assign when_LsuL1Plugin_l381 = LsuL1Plugin_logic_refill_free[0];
  assign when_LsuL1Plugin_l377_1 = (LsuL1Plugin_logic_refill_push_valid && LsuL1Plugin_logic_refill_free[1]);
  assign when_LsuL1Plugin_l381_1 = LsuL1Plugin_logic_refill_free[1];
  assign LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_refill_slots_0_valid && (! LsuL1Plugin_logic_refill_slots_0_cmdSent)) && (LsuL1Plugin_logic_refill_slots_0_victim == 2'b00));
  assign LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_1_0 = ((LsuL1Plugin_logic_refill_slots_1_valid && (! LsuL1Plugin_logic_refill_slots_1_cmdSent)) && (LsuL1Plugin_logic_refill_slots_1_victim == 2'b00));
  assign LsuL1Plugin_logic_refill_read_arbiter_hits = {LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_1_0,LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0};
  assign LsuL1Plugin_logic_refill_read_arbiter_hit = (|LsuL1Plugin_logic_refill_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_arbiter_oh = (LsuL1Plugin_logic_refill_read_arbiter_hits & {((LsuL1Plugin_logic_refill_read_arbiter_hits[0] & LsuL1Plugin_logic_refill_slots_1_priority) == 1'b0),((LsuL1Plugin_logic_refill_read_arbiter_hits[1] & LsuL1Plugin_logic_refill_slots_0_priority) == 1'b0)});
    if(when_LsuL1Plugin_l301) begin
      LsuL1Plugin_logic_refill_read_arbiter_oh = LsuL1Plugin_logic_refill_read_arbiter_lock;
    end
  end

  assign _zz_LsuL1Plugin_logic_refill_read_arbiter_sel = LsuL1Plugin_logic_refill_read_arbiter_oh[1];
  assign LsuL1Plugin_logic_refill_read_arbiter_sel = _zz_LsuL1Plugin_logic_refill_read_arbiter_sel;
  assign when_LsuL1Plugin_l301 = (|LsuL1Plugin_logic_refill_read_arbiter_lock);
  assign LsuL1Plugin_logic_bus_read_cmd_fire = (LsuL1Plugin_logic_bus_read_cmd_valid && LsuL1Plugin_logic_bus_read_cmd_ready);
  assign LsuL1Plugin_logic_refill_read_cmdAddress = {_zz_LsuL1Plugin_logic_refill_read_cmdAddress,6'h0};
  assign LsuL1Plugin_logic_bus_read_cmd_valid = LsuL1Plugin_logic_refill_read_arbiter_hit;
  assign LsuL1Plugin_logic_bus_read_cmd_payload_id = LsuL1Plugin_logic_refill_read_arbiter_sel;
  assign LsuL1Plugin_logic_bus_read_cmd_payload_address = LsuL1Plugin_logic_refill_read_cmdAddress;
  assign LsuL1Plugin_logic_refill_read_rspAddress = _zz_LsuL1Plugin_logic_refill_read_rspAddress;
  assign LsuL1Plugin_logic_refill_read_dirty = _zz_LsuL1Plugin_logic_refill_read_dirty;
  assign LsuL1Plugin_logic_refill_read_way = _zz_LsuL1Plugin_logic_refill_read_way;
  assign LsuL1Plugin_logic_refill_read_rspWithData = 1'b1;
  always @(*) begin
    LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_bankWriteNotif[0] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b0));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[1] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b1));
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_mask[0] = LsuL1Plugin_logic_refill_read_bankWriteNotif[0];
    LsuL1Plugin_logic_banksWrite_mask[1] = LsuL1Plugin_logic_refill_read_bankWriteNotif[1];
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      if(when_LsuL1Plugin_l929) begin
        LsuL1Plugin_logic_banksWrite_mask[0] = ((1'b0 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l929_1) begin
        LsuL1Plugin_logic_banksWrite_mask[1] = ((1'b1 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
    end
  end

  assign when_LsuL1Plugin_l450 = (LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_reservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_read_faulty = (LsuL1Plugin_logic_refill_read_hadError || LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refillCompletions = 2'b00;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refillCompletions[LsuL1Plugin_logic_bus_read_rsp_payload_id] = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_bus_read_rsp_ready = 1'b1;
  assign when_LsuL1Plugin_l463 = ((LsuL1Plugin_logic_refill_read_wordIndex == 1'b1) || (! LsuL1Plugin_logic_refill_read_rspWithData));
  assign LsuL1_REFILL_BUSY = {((! LsuL1Plugin_logic_refill_slots_1_loaded) && (! LsuL1Plugin_logic_refill_slots_1_loadedSet)),((! LsuL1Plugin_logic_refill_slots_0_loaded) && (! LsuL1Plugin_logic_refill_slots_0_loadedSet))};
  always @(*) begin
    LsuL1Plugin_logic_writeback_slots_0_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_write_rsp_valid) begin
      case(LsuL1Plugin_logic_bus_write_rsp_payload_id)
        1'b0 : begin
          LsuL1Plugin_logic_writeback_slots_0_fire = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign LsuL1Plugin_logic_writeback_slots_0_timer_done = (LsuL1Plugin_logic_writeback_slots_0_timer_counter == 1'b1);
  assign when_LsuL1Plugin_l530 = (LsuL1Plugin_logic_writeback_slots_0_timer_done && (LsuL1Plugin_logic_writeback_slots_0_fire || (! LsuL1Plugin_logic_writeback_slots_0_busy)));
  assign LsuL1Plugin_logic_writeback_slots_0_free = (! LsuL1Plugin_logic_writeback_slots_0_valid);
  always @(*) begin
    LsuL1Plugin_logic_writeback_slots_1_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_write_rsp_valid) begin
      case(LsuL1Plugin_logic_bus_write_rsp_payload_id)
        1'b0 : begin
        end
        default : begin
          LsuL1Plugin_logic_writeback_slots_1_fire = 1'b1;
        end
      endcase
    end
  end

  assign LsuL1Plugin_logic_writeback_slots_1_timer_done = (LsuL1Plugin_logic_writeback_slots_1_timer_counter == 1'b1);
  assign when_LsuL1Plugin_l530_1 = (LsuL1Plugin_logic_writeback_slots_1_timer_done && (LsuL1Plugin_logic_writeback_slots_1_fire || (! LsuL1Plugin_logic_writeback_slots_1_busy)));
  assign LsuL1Plugin_logic_writeback_slots_1_free = (! LsuL1Plugin_logic_writeback_slots_1_valid);
  assign LsuL1_WRITEBACK_BUSY = {(LsuL1Plugin_logic_writeback_slots_1_valid || LsuL1Plugin_logic_writeback_slots_1_fire),(LsuL1Plugin_logic_writeback_slots_0_valid || LsuL1Plugin_logic_writeback_slots_0_fire)};
  assign LsuL1Plugin_logic_writebackBusy = (|{LsuL1Plugin_logic_writeback_slots_1_valid,LsuL1Plugin_logic_writeback_slots_0_valid});
  assign _zz_LsuL1Plugin_logic_writeback_free = {LsuL1Plugin_logic_writeback_slots_1_free,LsuL1Plugin_logic_writeback_slots_0_free};
  assign LsuL1Plugin_logic_writeback_free = {_zz_LsuL1Plugin_logic_writeback_free_1[1],LsuL1Plugin_logic_writeback_slots_0_free};
  assign LsuL1Plugin_logic_writeback_full = (&{(! LsuL1Plugin_logic_writeback_slots_1_free),(! LsuL1Plugin_logic_writeback_slots_0_free)});
  always @(*) begin
    LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_valid = LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_waysWrite_tag_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_writeback_push_payload_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_way = 1'bx;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign when_LsuL1Plugin_l556 = (LsuL1Plugin_logic_writeback_free[0] && LsuL1Plugin_logic_writeback_push_valid);
  assign when_LsuL1Plugin_l561 = LsuL1Plugin_logic_writeback_free[0];
  assign when_LsuL1Plugin_l556_1 = (LsuL1Plugin_logic_writeback_free[1] && LsuL1Plugin_logic_writeback_push_valid);
  assign when_LsuL1Plugin_l561_1 = LsuL1Plugin_logic_writeback_free[1];
  assign LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0 = (LsuL1Plugin_logic_writeback_slots_0_valid && (! LsuL1Plugin_logic_writeback_slots_0_readCmdDone));
  assign LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_1_0 = (LsuL1Plugin_logic_writeback_slots_1_valid && (! LsuL1Plugin_logic_writeback_slots_1_readCmdDone));
  assign LsuL1Plugin_logic_writeback_read_arbiter_hits = {LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_1_0,LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0};
  assign LsuL1Plugin_logic_writeback_read_arbiter_hit = (|LsuL1Plugin_logic_writeback_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_read_arbiter_oh = (LsuL1Plugin_logic_writeback_read_arbiter_hits & {((LsuL1Plugin_logic_writeback_read_arbiter_hits[0] & LsuL1Plugin_logic_writeback_slots_1_priority) == 1'b0),((LsuL1Plugin_logic_writeback_read_arbiter_hits[1] & LsuL1Plugin_logic_writeback_slots_0_priority) == 1'b0)});
    if(when_LsuL1Plugin_l301_1) begin
      LsuL1Plugin_logic_writeback_read_arbiter_oh = LsuL1Plugin_logic_writeback_read_arbiter_lock;
    end
  end

  assign _zz_LsuL1Plugin_logic_writeback_read_arbiter_sel = LsuL1Plugin_logic_writeback_read_arbiter_oh[1];
  assign LsuL1Plugin_logic_writeback_read_arbiter_sel = _zz_LsuL1Plugin_logic_writeback_read_arbiter_sel;
  assign when_LsuL1Plugin_l301_1 = (|LsuL1Plugin_logic_writeback_read_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_read_address = _zz_LsuL1Plugin_logic_writeback_read_address;
  assign LsuL1Plugin_logic_writeback_read_way = _zz_LsuL1Plugin_logic_writeback_read_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_valid = LsuL1Plugin_logic_writeback_read_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_id = LsuL1Plugin_logic_writeback_read_arbiter_sel;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex = LsuL1Plugin_logic_writeback_read_wordIndex;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_way = LsuL1Plugin_logic_writeback_read_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_last = (LsuL1Plugin_logic_writeback_read_wordIndex == 1'b1);
  assign when_LsuL1Plugin_l605 = (LsuL1Plugin_logic_writeback_read_slotRead_valid && LsuL1Plugin_logic_writeback_read_slotRead_payload_last);
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_valid = LsuL1Plugin_logic_banks_0_usedByWriteback;
    if(when_LsuL1Plugin_l718) begin
      LsuL1Plugin_logic_banks_0_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_0_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b0));
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719) begin
      LsuL1Plugin_logic_banks_0_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_valid = LsuL1Plugin_logic_banks_1_usedByWriteback;
    if(when_LsuL1Plugin_l718_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_1_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b1));
  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  assign LsuL1Plugin_logic_writeback_read_readedData = _zz_LsuL1Plugin_logic_writeback_read_readedData;
  assign LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_writeback_slots_0_valid && LsuL1Plugin_logic_writeback_slots_0_victimBufferReady) && (! LsuL1Plugin_logic_writeback_slots_0_writeCmdDone));
  assign LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_1_0 = ((LsuL1Plugin_logic_writeback_slots_1_valid && LsuL1Plugin_logic_writeback_slots_1_victimBufferReady) && (! LsuL1Plugin_logic_writeback_slots_1_writeCmdDone));
  assign LsuL1Plugin_logic_writeback_write_arbiter_hits = {LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_1_0,LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0};
  assign LsuL1Plugin_logic_writeback_write_arbiter_hit = (|LsuL1Plugin_logic_writeback_write_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_arbiter_oh = (LsuL1Plugin_logic_writeback_write_arbiter_hits & {((LsuL1Plugin_logic_writeback_write_arbiter_hits[0] & LsuL1Plugin_logic_writeback_slots_1_priority) == 1'b0),((LsuL1Plugin_logic_writeback_write_arbiter_hits[1] & LsuL1Plugin_logic_writeback_slots_0_priority) == 1'b0)});
    if(when_LsuL1Plugin_l301_2) begin
      LsuL1Plugin_logic_writeback_write_arbiter_oh = LsuL1Plugin_logic_writeback_write_arbiter_lock;
    end
  end

  assign _zz_LsuL1Plugin_logic_writeback_write_arbiter_sel = LsuL1Plugin_logic_writeback_write_arbiter_oh[1];
  assign LsuL1Plugin_logic_writeback_write_arbiter_sel = _zz_LsuL1Plugin_logic_writeback_write_arbiter_sel;
  assign when_LsuL1Plugin_l301_2 = (|LsuL1Plugin_logic_writeback_write_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_write_last = (LsuL1Plugin_logic_writeback_write_wordIndex == 1'b1);
  assign LsuL1Plugin_logic_writeback_write_bufferRead_valid = LsuL1Plugin_logic_writeback_write_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_id = LsuL1Plugin_logic_writeback_write_arbiter_sel;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_last = LsuL1Plugin_logic_writeback_write_last;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = _zz_LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_fire = (LsuL1Plugin_logic_writeback_write_bufferRead_valid && LsuL1Plugin_logic_writeback_write_bufferRead_ready);
  assign when_LsuL1Plugin_l676 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && LsuL1Plugin_logic_writeback_write_last);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_bufferRead_ready = LsuL1Plugin_logic_writeback_write_cmd_ready;
    if(when_Stream_l477) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! LsuL1Plugin_logic_writeback_write_cmd_valid);
  assign LsuL1Plugin_logic_writeback_write_cmd_valid = LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_id = LsuL1Plugin_logic_writeback_write_bufferRead_rData_id;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_address = LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  assign _zz_LsuL1Plugin_logic_writeback_write_word = {LsuL1Plugin_logic_writeback_write_bufferRead_payload_id,LsuL1Plugin_logic_writeback_write_wordIndex};
  assign LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  assign LsuL1Plugin_logic_bus_write_cmd_valid = LsuL1Plugin_logic_writeback_write_cmd_valid;
  assign LsuL1Plugin_logic_writeback_write_cmd_ready = LsuL1Plugin_logic_bus_write_cmd_ready;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address = LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data = LsuL1Plugin_logic_writeback_write_word;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_id = LsuL1Plugin_logic_writeback_write_cmd_payload_id;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  assign LsuL1Plugin_logic_lsu_rb0_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 5];
  always @(*) begin
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[0] = LsuL1Plugin_logic_banks_0_usedByWriteback;
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1] = LsuL1Plugin_logic_banks_1_usedByWriteback;
  end

  assign when_LsuL1Plugin_l718 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719 = (! LsuL1Plugin_logic_banks_0_usedByWriteback);
  assign when_LsuL1Plugin_l718_1 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719_1 = (! LsuL1Plugin_logic_banks_1_usedByWriteback);
  assign when_LsuL1Plugin_l735 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0 = LsuL1Plugin_logic_banks_0_read_rsp;
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b0] || LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg);
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b1] || LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg);
  end

  assign when_LsuL1Plugin_l735_1 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1 = LsuL1Plugin_logic_banks_1_read_rsp;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 : 64'h0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 : 64'h0));
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0] = ((execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 3] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 3])) && 1'b1);
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1] = ((execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 3] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 3])) && 1'b1);
  end

  assign LsuL1Plugin_logic_shared_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_shared_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = LsuL1Plugin_logic_shared_write_payload_data_dirty;
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
    end
  end

  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = LsuL1Plugin_logic_shared_lsuRead_rsp_dirty;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = LsuL1Plugin_logic_ways_0_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = LsuL1Plugin_logic_ways_1_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault;
  assign LsuL1Plugin_logic_lsu_sharedBypassers_0_hit = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0 = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_plru_0 : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0);
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_dirty : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty);
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
  end

  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 = (|execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0);
  assign execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0 = (execute_ctrl4_down_LsuL1_STORE_lane0 || execute_ctrl4_down_LsuL1_ATOMIC_lane0);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0 = (! LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0[0] = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id[0];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0 = execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazards = {(LsuL1Plugin_logic_refill_slots_1_valid && (LsuL1Plugin_logic_refill_slots_1_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6])),(LsuL1Plugin_logic_refill_slots_0_valid && (LsuL1Plugin_logic_refill_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]))};
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazards = {(LsuL1Plugin_logic_writeback_slots_1_valid && (LsuL1Plugin_logic_writeback_slots_1_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6])),(LsuL1Plugin_logic_writeback_slots_0_valid && (LsuL1Plugin_logic_writeback_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]))};
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazard = (|LsuL1Plugin_logic_lsu_ctrl_refillHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazard = (|LsuL1Plugin_logic_lsu_ctrl_writebackHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_wasDirty = (|(execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadedDirties = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty = LsuL1Plugin_logic_lsu_ctrl_loadedDirties[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_bankNotRead = (|(execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadHazard = ((execute_ctrl4_down_LsuL1_LOAD_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (LsuL1Plugin_logic_lsu_ctrl_bankNotRead || LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_storeHazard = ((execute_ctrl4_down_LsuL1_STORE_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (! LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_preventSideEffects = (execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_freeze_valid);
  assign LsuL1Plugin_logic_lsu_ctrl_flushHazard = (execute_ctrl4_down_LsuL1_FLUSH_lane0 && (! LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_coherencyHazard = 1'b0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0 = 1'b0;
  assign execute_ctrl4_down_LsuL1_HAZARD_lane0 = (((((LsuL1Plugin_logic_lsu_ctrl_hazardReg || LsuL1Plugin_logic_lsu_ctrl_loadHazard) || LsuL1Plugin_logic_lsu_ctrl_refillHazard) || LsuL1Plugin_logic_lsu_ctrl_storeHazard) || LsuL1Plugin_logic_lsu_ctrl_coherencyHazard) || execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0);
  assign execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 = (LsuL1Plugin_logic_lsu_ctrl_flushHazardReg || LsuL1Plugin_logic_lsu_ctrl_flushHazard);
  assign execute_ctrl4_down_LsuL1_MISS_lane0 = (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0);
  assign execute_ctrl4_down_LsuL1_FAULT_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (|(execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 & {execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault}))) && (! execute_ctrl4_down_LsuL1_FLUSH_lane0));
  assign execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0) && 1'b0);
  assign execute_ctrl4_down_LsuL1_REFILL_HIT_lane0 = LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  assign LsuL1Plugin_logic_lsu_ctrl_canRefill = (((! (LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_refill_full)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_canFlush = (((LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win && (! LsuL1Plugin_logic_writeback_full)) && (! (|{LsuL1Plugin_logic_refill_slots_1_valid,LsuL1Plugin_logic_refill_slots_0_valid}))) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs = LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[1];
  always @(*) begin
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[0] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 && (! LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0));
  end

  assign LsuL1Plugin_logic_lsu_ctrl_needFlushOh = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel = LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushSel = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  assign LsuL1Plugin_logic_lsu_ctrl_isAccess = (((! execute_ctrl4_down_LsuL1_FLUSH_lane0) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_askRefill = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askUpgrade = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askFlush = ((execute_ctrl4_down_LsuL1_FLUSH_lane0 && LsuL1Plugin_logic_lsu_ctrl_canFlush) && (|LsuL1Plugin_logic_lsu_ctrl_needFlushs));
  assign LsuL1Plugin_logic_lsu_ctrl_askCbm = (execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (execute_ctrl4_down_LsuL1_INVALID_lane0 || (execute_ctrl4_down_LsuL1_CLEAN_lane0 && LsuL1Plugin_logic_lsu_ctrl_wasDirty)));
  assign LsuL1Plugin_logic_lsu_ctrl_doRefill = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_doUpgrade = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askUpgrade);
  assign LsuL1Plugin_logic_lsu_ctrl_doFlush = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askFlush);
  assign LsuL1Plugin_logic_lsu_ctrl_doWrite = ((((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_STORE_lane0) && execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0) && _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite[0]) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_doCbm = (((((execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askCbm) && LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) && (! LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_lsu_ctrl_refillHazard)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_wayId = _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  assign LsuL1Plugin_logic_lsu_ctrl_targetWay = (LsuL1Plugin_logic_lsu_ctrl_askUpgrade ? LsuL1Plugin_logic_lsu_ctrl_wayId : LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_wayId;
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_doRefillPush = (LsuL1Plugin_logic_lsu_ctrl_doRefill || LsuL1Plugin_logic_lsu_ctrl_doUpgrade);
  always @(*) begin
    LsuL1Plugin_logic_refill_push_valid = LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_refill_push_valid = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_unique = execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_data = LsuL1Plugin_logic_lsu_ctrl_askRefill;
  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_wayId;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_victim = ((LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty) ? LsuL1Plugin_logic_writeback_free : 2'b00);
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_victim = 2'b00;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_dirty = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0 = (LsuL1Plugin_logic_lsu_ctrl_refillHazards | (((! execute_ctrl4_down_LsuL1_HAZARD_lane0) && (LsuL1Plugin_logic_lsu_ctrl_askRefill || LsuL1Plugin_logic_lsu_ctrl_askUpgrade)) ? (LsuL1Plugin_logic_refill_full ? 2'b11 : LsuL1Plugin_logic_refill_free) : 2'b00));
  assign execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0 = 2'b00;
  assign when_LsuL1Plugin_l915 = (execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_ABORD_lane0));
  assign _zz_23 = {LsuL1Plugin_logic_lsu_ctrl_askRefill,{LsuL1Plugin_logic_lsu_ctrl_doUpgrade,LsuL1Plugin_logic_lsu_ctrl_doFlush}};
  always @(*) begin
    LsuL1Plugin_logic_shared_write_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(when_LsuL1Plugin_l1018) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b0;
    end
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_shared_write_payload_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_plru_0 = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_shared_write_payload_data_plru_0 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1[0 : 0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_dirty = ((execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty | (LsuL1Plugin_logic_lsu_ctrl_doWrite ? execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 : 2'b00)) & (~ ((LsuL1Plugin_logic_lsu_ctrl_doRefill ? _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty : 2'b00) | (LsuL1Plugin_logic_lsu_ctrl_doFlush ? LsuL1Plugin_logic_lsu_ctrl_needFlushOh : 2'b00))));
    if(when_LsuL1Plugin_l1218) begin
      LsuL1Plugin_logic_shared_write_payload_data_dirty = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[2 : 1];
    end
  end

  assign _zz_24 = ({3'd0,1'b1} <<< execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[4 : 3]);
  assign when_LsuL1Plugin_l929 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign when_LsuL1Plugin_l929_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 = (|LsuL1Plugin_logic_lsu_ctrl_needFlushs);
  assign _zz_LsuL1Plugin_logic_waysWrite_tag_address = _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = LsuL1Plugin_logic_lsu_ctrl_doWrite;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign when_LsuL1Plugin_l1018 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0));
  always @(*) begin
    execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
    if(when_LsuL1Plugin_l1025) begin
      if(when_LsuL1Plugin_l1029) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1029_1) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1029_2) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1029_3) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
      if(when_LsuL1Plugin_l1029_4) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[39 : 32] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[39 : 32];
      end
      if(when_LsuL1Plugin_l1029_5) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[47 : 40] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[47 : 40];
      end
      if(when_LsuL1Plugin_l1029_6) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[55 : 48] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[55 : 48];
      end
      if(when_LsuL1Plugin_l1029_7) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[63 : 56] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[63 : 56];
      end
    end
    if(when_LsuL1Plugin_l1025_1) begin
      if(when_LsuL1Plugin_l1029_8) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1029_9) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1029_10) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1029_11) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
      if(when_LsuL1Plugin_l1029_12) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[39 : 32] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[39 : 32];
      end
      if(when_LsuL1Plugin_l1029_13) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[47 : 40] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[47 : 40];
      end
      if(when_LsuL1Plugin_l1029_14) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[55 : 48] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[55 : 48];
      end
      if(when_LsuL1Plugin_l1029_15) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[63 : 56] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[63 : 56];
      end
    end
  end

  assign when_LsuL1Plugin_l1025 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1];
  assign when_LsuL1Plugin_l1029 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1029_1 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1029_2 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1029_3 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l1029_4 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[4];
  assign when_LsuL1Plugin_l1029_5 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[5];
  assign when_LsuL1Plugin_l1029_6 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[6];
  assign when_LsuL1Plugin_l1029_7 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[7];
  assign when_LsuL1Plugin_l1025_1 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0];
  assign when_LsuL1Plugin_l1029_8 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1029_9 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1029_10 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1029_11 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l1029_12 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[4];
  assign when_LsuL1Plugin_l1029_13 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[5];
  assign when_LsuL1Plugin_l1029_14 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[6];
  assign when_LsuL1Plugin_l1029_15 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[7];
  assign execute_ctrl4_down_LsuL1_READ_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  assign LsuL1Plugin_logic_initializer_done = LsuL1Plugin_logic_initializer_counter[6];
  assign when_LsuL1Plugin_l1218 = (! LsuL1Plugin_logic_initializer_done);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0 = 3'b000;
  assign LsuL1Plugin_logic_refill_read_reservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_reservation_take));
  assign LsuL1Plugin_logic_refill_read_writeReservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_writeReservation_take));
  assign PrefetcherRptPlugin_logic_order_ready = PrefetcherRptPlugin_logic_order_fifo_io_push_ready;
  assign PrefetcherRptPlugin_logic_queued_valid = PrefetcherRptPlugin_logic_order_fifo_io_pop_valid;
  assign PrefetcherRptPlugin_logic_queued_payload_address = PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_address;
  assign PrefetcherRptPlugin_logic_queued_payload_unique = PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_unique;
  assign PrefetcherRptPlugin_logic_queued_payload_from = PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_from;
  assign PrefetcherRptPlugin_logic_queued_payload_to = PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_to;
  assign PrefetcherRptPlugin_logic_queued_payload_stride = PrefetcherRptPlugin_logic_order_fifo_io_pop_payload_stride;
  assign PrefetcherRptPlugin_logic_advanceAt = (PrefetcherRptPlugin_logic_queued_payload_from + PrefetcherRptPlugin_logic_counter);
  assign PrefetcherRptPlugin_logic_done = (PrefetcherRptPlugin_logic_advanceAt == PrefetcherRptPlugin_logic_queued_payload_to);
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_valid = PrefetcherRptPlugin_logic_queued_valid;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_address = PrefetcherRptPlugin_logic_queued_payload_address;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_unique = PrefetcherRptPlugin_logic_queued_payload_unique;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_from = PrefetcherRptPlugin_logic_queued_payload_from;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_to = PrefetcherRptPlugin_logic_queued_payload_to;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_payload_stride = PrefetcherRptPlugin_logic_queued_payload_stride;
  assign PrefetcherRptPlugin_logic_queued_ready = (PrefetcherRptPlugin_logic_queued_forkSerial_next_ready && PrefetcherRptPlugin_logic_done);
  assign PrefetcherRptPlugin_logic_pip2_node_0_valid = PrefetcherRptPlugin_logic_queued_forkSerial_next_valid;
  assign PrefetcherRptPlugin_logic_queued_forkSerial_next_ready = (PrefetcherRptPlugin_logic_pip2_node_0_isReady || PrefetcherRptPlugin_logic_pip2_node_0_isCancel);
  assign PrefetcherRptPlugin_logic_pip2_node_0_CMD_address = PrefetcherRptPlugin_logic_queued_payload_address;
  assign PrefetcherRptPlugin_logic_pip2_node_0_CMD_unique = PrefetcherRptPlugin_logic_queued_payload_unique;
  assign PrefetcherRptPlugin_logic_pip2_node_0_CMD_from = PrefetcherRptPlugin_logic_queued_payload_from;
  assign PrefetcherRptPlugin_logic_pip2_node_0_CMD_to = PrefetcherRptPlugin_logic_queued_payload_to;
  assign PrefetcherRptPlugin_logic_pip2_node_0_CMD_stride = PrefetcherRptPlugin_logic_queued_payload_stride;
  assign PrefetcherRptPlugin_logic_pip2_node_0_MUL = ($signed(_zz_PrefetcherRptPlugin_logic_pip2_node_0_MUL) * $signed(PrefetcherRptPlugin_logic_queued_payload_stride));
  assign PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR = _zz_PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR;
  assign PrefetcherRptPlugin_io_valid = PrefetcherRptPlugin_logic_pip2_node_1_isValid;
  assign PrefetcherRptPlugin_logic_pip2_node_1_ready = PrefetcherRptPlugin_io_ready;
  assign PrefetcherRptPlugin_io_payload_address = PrefetcherRptPlugin_logic_pip2_node_1_adder_ADDR;
  assign PrefetcherRptPlugin_io_payload_unique = PrefetcherRptPlugin_logic_pip2_node_1_CMD_unique;
  always @(*) begin
    PrefetcherRptPlugin_logic_pip2_node_0_ready = PrefetcherRptPlugin_logic_pip2_node_1_ready;
    if(when_StageLink_l71) begin
      PrefetcherRptPlugin_logic_pip2_node_0_ready = 1'b1;
    end
  end

  assign when_StageLink_l71 = (! PrefetcherRptPlugin_logic_pip2_node_1_isValid);
  assign PrefetcherRptPlugin_logic_pip2_node_0_isFiring = (PrefetcherRptPlugin_logic_pip2_node_0_isValid && PrefetcherRptPlugin_logic_pip2_node_0_isReady);
  assign PrefetcherRptPlugin_logic_pip2_node_0_isValid = PrefetcherRptPlugin_logic_pip2_node_0_valid;
  assign PrefetcherRptPlugin_logic_pip2_node_0_isReady = PrefetcherRptPlugin_logic_pip2_node_0_ready;
  assign PrefetcherRptPlugin_logic_pip2_node_0_isCancel = 1'b0;
  assign PrefetcherRptPlugin_logic_pip2_node_1_isValid = PrefetcherRptPlugin_logic_pip2_node_1_valid;
  assign _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag = PrefetcherRptPlugin_logic_storage_ram_spinal_port0;
  assign PrefetcherRptPlugin_logic_storage_read_rsp_tag = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[14 : 0];
  assign PrefetcherRptPlugin_logic_storage_read_rsp_address = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[30 : 15];
  assign PrefetcherRptPlugin_logic_storage_read_rsp_stride = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[42 : 31];
  assign PrefetcherRptPlugin_logic_storage_read_rsp_score = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[47 : 43];
  assign PrefetcherRptPlugin_logic_storage_read_rsp_advance = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[50 : 48];
  assign PrefetcherRptPlugin_logic_storage_read_rsp_missed = _zz_PrefetcherRptPlugin_logic_storage_read_rsp_tag[51];
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0 = execute_ctrl2_up_integer_RS1_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 = execute_ctrl2_up_integer_RS2_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0[31]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0[31]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        if(when_TrapPlugin_l654) begin
          PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_harts_0_int_pending = 1'b0;
    if(TrapPlugin_logic_harts_0_interrupt_pendingInterrupt) begin
      PrivilegedPlugin_logic_harts_0_int_pending = 1'b1;
    end
  end

  assign PrivilegedPlugin_logic_harts_0_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_hartRunning = 1'b1;
  assign PrivilegedPlugin_logic_harts_0_debugMode = (! PrivilegedPlugin_logic_harts_0_hartRunning);
  assign PrivilegedPlugin_logic_harts_0_m_status_mpp = 2'b11;
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b0;
    if(when_PrivilegedPlugin_l554) begin
      PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b1;
    end
  end

  assign PrivilegedPlugin_logic_harts_0_m_status_tw = 1'b0;
  assign when_PrivilegedPlugin_l549 = (PrivilegedPlugin_logic_harts_0_m_status_fs != 2'b00);
  assign when_PrivilegedPlugin_l550 = (|FpuCsrPlugin_api_gotDirty);
  assign when_PrivilegedPlugin_l554 = (PrivilegedPlugin_logic_harts_0_m_status_fs == 2'b11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_768);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_834);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_836);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue && REG_CSR_772);
  assign _zz_when_TrapPlugin_l207 = (PrivilegedPlugin_logic_harts_0_m_ip_mtip && PrivilegedPlugin_logic_harts_0_m_ie_mtie);
  assign _zz_when_TrapPlugin_l207_1 = (PrivilegedPlugin_logic_harts_0_m_ip_msip && PrivilegedPlugin_logic_harts_0_m_ie_msie);
  assign _zz_when_TrapPlugin_l207_2 = (PrivilegedPlugin_logic_harts_0_m_ip_meip && PrivilegedPlugin_logic_harts_0_m_ie_meie);
  always @(*) begin
    case(execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 & execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 | execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 ^ execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        late0_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign late0_IntAluPlugin_logic_alu_result = (_zz_late0_IntAluPlugin_logic_alu_result | _zz_late0_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0 = late0_IntAluPlugin_logic_alu_result;
  assign late0_IntAluPlugin_logic_wb_valid = execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0;
  assign late0_IntAluPlugin_logic_wb_payload = execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0;
  assign late0_BarrelShifterPlugin_logic_shift_amplitude = _zz_late0_BarrelShifterPlugin_logic_shift_amplitude;
  assign late0_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_late0_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0);
  assign late0_BarrelShifterPlugin_logic_shift_shifted = _zz_late0_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign late0_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_late0_BarrelShifterPlugin_logic_shift_patched : late0_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = late0_BarrelShifterPlugin_logic_shift_patched;
  assign late0_BarrelShifterPlugin_logic_wb_valid = execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0;
  assign late0_BarrelShifterPlugin_logic_wb_payload = execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  always @(*) begin
    case(execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 & execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 | execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 ^ execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      default : begin
        early1_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign early1_IntAluPlugin_logic_alu_result = (_zz_early1_IntAluPlugin_logic_alu_result | _zz_early1_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1 = early1_IntAluPlugin_logic_alu_result;
  assign early1_IntAluPlugin_logic_wb_valid = execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1;
  assign early1_IntAluPlugin_logic_wb_payload = execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1;
  assign early1_BarrelShifterPlugin_logic_shift_amplitude = _zz_early1_BarrelShifterPlugin_logic_shift_amplitude;
  assign early1_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_early1_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1);
  assign early1_BarrelShifterPlugin_logic_shift_shifted = _zz_early1_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign early1_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_early1_BarrelShifterPlugin_logic_shift_patched : early1_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1 = early1_BarrelShifterPlugin_logic_shift_patched;
  assign early1_BarrelShifterPlugin_logic_wb_valid = execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1;
  assign early1_BarrelShifterPlugin_logic_wb_payload = execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  always @(*) begin
    case(execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 & execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 | execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 ^ execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      default : begin
        late1_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign late1_IntAluPlugin_logic_alu_result = (_zz_late1_IntAluPlugin_logic_alu_result | _zz_late1_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1 = late1_IntAluPlugin_logic_alu_result;
  assign late1_IntAluPlugin_logic_wb_valid = execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1;
  assign late1_IntAluPlugin_logic_wb_payload = execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1;
  assign late1_BarrelShifterPlugin_logic_shift_amplitude = _zz_late1_BarrelShifterPlugin_logic_shift_amplitude;
  assign late1_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_late1_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1);
  assign late1_BarrelShifterPlugin_logic_shift_shifted = _zz_late1_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign late1_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_late1_BarrelShifterPlugin_logic_shift_patched : late1_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1 = late1_BarrelShifterPlugin_logic_shift_patched;
  assign late1_BarrelShifterPlugin_logic_wb_valid = execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1;
  assign late1_BarrelShifterPlugin_logic_wb_payload = execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  assign FpuMvPlugin_logic_iwb_valid = execute_ctrl3_down_FpuMvPlugin_SEL_INT_lane0;
  assign FpuMvPlugin_logic_iwb_payload = execute_ctrl3_up_float_RS1_lane0[31:0];
  assign FpuMvPlugin_logic_fwb_valid = execute_ctrl4_down_FpuMvPlugin_SEL_FLOAT_lane0;
  always @(*) begin
    FpuMvPlugin_logic_fwb_payload[31 : 0] = execute_ctrl4_up_integer_RS1_lane0[31 : 0];
    FpuMvPlugin_logic_fwb_payload[63 : 32] = 32'hffffffff;
  end

  assign WhiteboxerPlugin_logic_fetch_fire = fetch_logic_ctrls_0_down_isFiring;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_valid = LsuL1Plugin_logic_bus_read_cmd_valid;
  assign LsuL1Plugin_logic_bus_read_cmd_ready = LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_ready;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_last = 1'b1;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_write = 1'b0;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_id = LsuL1Plugin_logic_bus_read_cmd_payload_id;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_payload_fragment_address = LsuL1Plugin_logic_bus_read_cmd_payload_address;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_valid = LsuL1Plugin_logic_bus_write_cmd_valid;
  assign LsuL1Plugin_logic_bus_write_cmd_ready = LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_ready;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_last = LsuL1Plugin_logic_bus_write_cmd_payload_last;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_write = 1'b1;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_id = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_id;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_payload_fragment_address = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_readCmd_ready = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_0_ready;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_writeCmd_ready = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_inputs_1_ready;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_fire = (LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_valid && LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready);
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_ready = (LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready && (LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_last == LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_last));
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_valid = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_valid;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_write = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_write;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_id = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_id;
  always @(*) begin
    LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_address = LsuL1Plugin_logic_bus_toWishbone_arbiter_arbiter_io_output_payload_fragment_address;
    LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_address[5 : 5] = LsuL1Plugin_logic_bus_toWishbone_arbiter_counter;
  end

  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_data = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_last = (&LsuL1Plugin_logic_bus_toWishbone_arbiter_counter);
  always @(*) begin
    LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_ready;
    if(when_Stream_l477_1) begin
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready = 1'b1;
    end
  end

  assign when_Stream_l477_1 = (! LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid);
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rValid;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_last = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_last;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_write = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_write;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_id = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_id;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_address = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_address;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_data = LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_data;
  assign LsuL1WishbonePlugin_logic_bus_ADR = (LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_address >>> 3'd5);
  assign LsuL1WishbonePlugin_logic_bus_CTI = (LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_last ? 3'b111 : 3'b010);
  assign LsuL1WishbonePlugin_logic_bus_BTE = 2'b00;
  assign LsuL1WishbonePlugin_logic_bus_SEL = 32'hffffffff;
  assign LsuL1WishbonePlugin_logic_bus_WE = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_write;
  assign LsuL1WishbonePlugin_logic_bus_DAT_MOSI = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_data;
  assign LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_ready = (LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid && (LsuL1WishbonePlugin_logic_bus_ACK || LsuL1WishbonePlugin_logic_bus_ERR));
  assign LsuL1WishbonePlugin_logic_bus_CYC = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid;
  assign LsuL1WishbonePlugin_logic_bus_STB = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid;
  assign LsuL1Plugin_logic_bus_read_rsp_valid = ((LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid && (! LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_write)) && (LsuL1WishbonePlugin_logic_bus_ACK || LsuL1WishbonePlugin_logic_bus_ERR));
  assign LsuL1Plugin_logic_bus_read_rsp_payload_error = LsuL1WishbonePlugin_logic_bus_ERR;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_id = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_id;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_data = LsuL1WishbonePlugin_logic_bus_DAT_MISO;
  assign LsuL1Plugin_logic_bus_write_rsp_valid = (((LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_valid && LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_write) && LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_last) && (LsuL1WishbonePlugin_logic_bus_ACK || LsuL1WishbonePlugin_logic_bus_ERR));
  assign LsuL1Plugin_logic_bus_write_rsp_payload_error = LsuL1WishbonePlugin_logic_bus_ERR;
  assign LsuL1Plugin_logic_bus_write_rsp_payload_id = LsuL1Plugin_logic_bus_toWishbone_arbiter_buffered_payload_fragment_id;
  always @(*) begin
    CsrAccessPlugin_bus_decode_exception = 1'b0;
    if(when_PrivilegedPlugin_l701) begin
      CsrAccessPlugin_bus_decode_exception = 1'b1;
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trap = 1'b0;
    if(when_CsrAccessPlugin_l155) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trapCode = 4'bxxxx;
    if(when_CsrAccessPlugin_l155) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_read_halt = 1'b0;
    if(when_CsrRamPlugin_l85) begin
      CsrAccessPlugin_bus_read_halt = 1'b1;
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_write_halt = 1'b0;
    if(when_CsrRamPlugin_l96) begin
      CsrAccessPlugin_bus_write_halt = 1'b1;
    end
  end

  assign FetchL1Plugin_logic_banks_0_read_rsp = FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0 = FetchL1Plugin_logic_banks_0_read_rsp;
  assign FetchL1Plugin_logic_banks_1_read_rsp = FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1 = FetchL1Plugin_logic_banks_1_read_rsp;
  always @(*) begin
    FetchL1Plugin_logic_waysWrite_mask = 2'b00;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_mask = 2'b11;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      if(when_FetchL1Plugin_l304) begin
        FetchL1Plugin_logic_waysWrite_mask[FetchL1Plugin_logic_refill_onRsp_wayToAllocate] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_refill_onRsp_address[11 : 6];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_error = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_address = FetchL1Plugin_logic_refill_onRsp_address[31 : 12];
    end
  end

  assign _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded = FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_0_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_0_read_rsp_error = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_0_read_rsp_address = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = FetchL1Plugin_logic_ways_0_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = FetchL1Plugin_logic_ways_0_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded = FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_1_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_1_read_rsp_error = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_1_read_rsp_address = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = FetchL1Plugin_logic_ways_1_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = FetchL1Plugin_logic_ways_1_read_rsp_address;
  assign FetchL1Plugin_logic_plru_read_rsp_0 = FetchL1Plugin_logic_plru_mem_spinal_port1[0 : 0];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0 = FetchL1Plugin_logic_plru_read_rsp_0;
  assign FetchL1Plugin_logic_invalidate_cmd_valid = (|TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid);
  always @(*) begin
    FetchL1Plugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchL1Plugin_l268) begin
      FetchL1Plugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_invalidate_counterIncr = (FetchL1Plugin_logic_invalidate_counter + 7'h01);
  assign FetchL1Plugin_logic_invalidate_done = FetchL1Plugin_logic_invalidate_counter[6];
  assign FetchL1Plugin_logic_invalidate_last = FetchL1Plugin_logic_invalidate_counterIncr[6];
  assign when_FetchL1Plugin_l204 = (! FetchL1Plugin_logic_invalidate_done);
  assign when_FetchL1Plugin_l211 = ((FetchL1Plugin_logic_invalidate_done && FetchL1Plugin_logic_invalidate_cmd_valid) && FetchL1Plugin_logic_invalidate_canStart);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      if(FetchL1Plugin_logic_invalidate_last) begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b1;
      end
    end
  end

  assign when_FetchL1Plugin_l216 = (! FetchL1Plugin_logic_invalidate_done);
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  assign FetchL1Plugin_logic_refill_slots_0_askCmd = (FetchL1Plugin_logic_refill_slots_0_valid && (! FetchL1Plugin_logic_refill_slots_0_cmdSent));
  assign FetchL1Plugin_logic_refill_slots_1_askCmd = (FetchL1Plugin_logic_refill_slots_1_valid && (! FetchL1Plugin_logic_refill_slots_1_cmdSent));
  assign when_FetchL1Plugin_l246 = (! FetchL1Plugin_logic_refill_slots_1_valid);
  assign when_FetchL1Plugin_l246_1 = (! FetchL1Plugin_logic_refill_slots_0_valid);
  assign _zz_38 = (! FetchL1Plugin_logic_refill_slots_0_valid);
  assign _zz_39 = {(! FetchL1Plugin_logic_refill_slots_1_valid),_zz_38};
  assign FetchL1Plugin_logic_refill_hazard = (|{(FetchL1Plugin_logic_refill_slots_1_valid && (FetchL1Plugin_logic_refill_slots_1_address[11 : 6] == FetchL1Plugin_logic_refill_start_address[11 : 6])),(FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == FetchL1Plugin_logic_refill_start_address[11 : 6]))});
  assign when_FetchL1Plugin_l255 = ((FetchL1Plugin_logic_refill_start_valid && FetchL1Plugin_logic_invalidate_done) && (! FetchL1Plugin_logic_refill_hazard));
  assign when_FetchL1Plugin_l268 = ((|{FetchL1Plugin_logic_refill_slots_1_valid,FetchL1Plugin_logic_refill_slots_0_valid}) || FetchL1Plugin_logic_refill_start_valid);
  assign FetchL1Plugin_logic_refill_onCmd_propoedOh = {(FetchL1Plugin_logic_refill_slots_1_askCmd && (&((! FetchL1Plugin_logic_refill_slots_0_askCmd) || (! FetchL1Plugin_logic_refill_slots_0_priority[1])))),(FetchL1Plugin_logic_refill_slots_0_askCmd && (&((! FetchL1Plugin_logic_refill_slots_1_askCmd) || (! FetchL1Plugin_logic_refill_slots_1_priority[0]))))};
  assign when_FetchL1Plugin_l276 = (! FetchL1Plugin_logic_refill_onCmd_locked);
  assign FetchL1Plugin_logic_refill_onCmd_oh = (FetchL1Plugin_logic_refill_onCmd_locked ? FetchL1Plugin_logic_refill_onCmd_lockedOh : FetchL1Plugin_logic_refill_onCmd_propoedOh);
  assign _zz_FetchL1Plugin_logic_bus_cmd_payload_address = FetchL1Plugin_logic_refill_onCmd_oh[0];
  assign _zz_FetchL1Plugin_logic_bus_cmd_payload_id = FetchL1Plugin_logic_refill_onCmd_oh[1];
  assign FetchL1Plugin_logic_bus_cmd_valid = (|FetchL1Plugin_logic_refill_onCmd_oh);
  assign FetchL1Plugin_logic_bus_cmd_payload_address = {((_zz_FetchL1Plugin_logic_bus_cmd_payload_address ? FetchL1Plugin_logic_refill_slots_0_address[31 : 6] : 26'h0) | (_zz_FetchL1Plugin_logic_bus_cmd_payload_id ? FetchL1Plugin_logic_refill_slots_1_address[31 : 6] : 26'h0)),6'h0};
  assign FetchL1Plugin_logic_bus_cmd_payload_io = _zz_FetchL1Plugin_logic_bus_cmd_payload_io[0];
  assign FetchL1Plugin_logic_bus_cmd_payload_id = _zz_FetchL1Plugin_logic_bus_cmd_payload_id;
  assign FetchL1Plugin_logic_refill_onRsp_holdHarts = ((|FetchL1Plugin_logic_waysWrite_mask) || (|{((FetchL1Plugin_logic_refill_slots_1_valid && (FetchL1Plugin_logic_refill_slots_1_address[11 : 6] == fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6])) && (! ((FetchL1Plugin_logic_refill_onRsp_rspIdReg == _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts) && (_zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_1 < FetchL1Plugin_logic_refill_onRsp_wordIndex)))),((FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6])) && (! ((FetchL1Plugin_logic_refill_onRsp_rspIdReg == _zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_2) && (_zz_FetchL1Plugin_logic_refill_onRsp_holdHarts_3 < FetchL1Plugin_logic_refill_onRsp_wordIndex))))}));
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297 = FetchL1Plugin_logic_refill_onRsp_holdHarts;
  assign FetchL1Plugin_logic_bus_rsp_fire = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_ready);
  assign FetchL1Plugin_logic_refill_onRsp_wayToAllocate = _zz_FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  assign FetchL1Plugin_logic_refill_onRsp_address = _zz_FetchL1Plugin_logic_refill_onRsp_address;
  assign when_FetchL1Plugin_l304 = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_firstCycle || FetchL1Plugin_logic_bus_rsp_payload_error));
  assign FetchL1Plugin_logic_banks_0_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b0));
  assign FetchL1Plugin_logic_banks_0_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_0_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_banks_1_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b1));
  assign FetchL1Plugin_logic_banks_1_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_1_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_ready = 1'b1;
  assign when_FetchL1Plugin_l330 = (FetchL1Plugin_logic_refill_onRsp_wordIndex == 1'b1);
  assign FetchL1Plugin_logic_cmd_doIt = (fetch_logic_ctrls_1_up_ready || ((! fetch_logic_ctrls_1_up_valid) && 1'b1));
  assign FetchL1Plugin_logic_banks_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 5];
  assign FetchL1Plugin_logic_banks_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 5];
  assign FetchL1Plugin_logic_ways_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_plru_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_plru_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = (FetchL1Plugin_logic_plru_write_valid && (FetchL1Plugin_logic_plru_write_payload_address == FetchL1Plugin_logic_plru_read_cmd_payload));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = FetchL1Plugin_logic_plru_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = (|FetchL1Plugin_logic_waysWrite_mask);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = FetchL1Plugin_logic_waysWrite_address;
  always @(*) begin
    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
    if(fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID) begin
      fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
    end
  end

  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_Fetch_WORD = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 : 64'h0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 : 64'h0));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS == fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 6]));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0 = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1 = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_TRANSLATED[31 : 12]));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT = (|{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1,fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0});
  assign FetchL1Plugin_logic_ctrl_pmaPort_cmd_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0 = (! FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id = FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0[0] = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0 = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  always @(*) begin
    FetchL1Plugin_logic_plru_write_valid = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_data_0 = _zz_FetchL1Plugin_logic_plru_write_payload_data_0[0 : 0];
    end
  end

  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isReady);
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address = fetch_logic_ctrls_2_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  assign FetchL1Plugin_logic_refill_start_wayToAllocate = FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  assign FetchL1Plugin_logic_ctrl_dataAccessFault = (_zz_FetchL1Plugin_logic_ctrl_dataAccessFault[0] && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
  always @(*) begin
    FetchL1Plugin_logic_trapPort_valid = 1'b0;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l533) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_trapPort_payload_tval = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_exception = 1'bx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_code = 4'bxxxx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
      if(when_FetchL1Plugin_l520) begin
        FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
      end
    end
  end

  assign _zz_71 = zz_FetchL1Plugin_logic_trapPort_payload_arg(1'b0);
  always @(*) FetchL1Plugin_logic_trapPort_payload_arg = _zz_71;
  always @(*) begin
    FetchL1Plugin_logic_ctrl_allowRefill = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
  end

  assign when_FetchL1Plugin_l474 = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD);
  assign when_FetchL1Plugin_l480 = ((FetchL1Plugin_logic_ctrl_dataAccessFault || FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT);
  assign when_FetchL1Plugin_l487 = (fetch_logic_ctrls_2_down_MMU_PAGE_FAULT || (! fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE));
  assign when_FetchL1Plugin_l520 = (! fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION);
  always @(*) begin
    FetchL1Plugin_logic_refill_start_valid = (FetchL1Plugin_logic_ctrl_allowRefill && (! FetchL1Plugin_logic_ctrl_trapSent));
    if(when_FetchL1Plugin_l537) begin
      FetchL1Plugin_logic_refill_start_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_refill_start_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_refill_start_isIo = FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  assign fetch_logic_ctrls_2_down_TRAP = (FetchL1Plugin_logic_trapPort_valid || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l533 = ((! fetch_logic_ctrls_2_up_isValid) || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l537 = ((! fetch_logic_ctrls_2_up_isValid) && 1'b1);
  assign when_FetchL1Plugin_l541 = (((! fetch_logic_ctrls_2_up_isValid) || fetch_logic_ctrls_2_down_isReady) || fetch_logic_ctrls_2_up_isCanceling);
  assign when_FetchL1Plugin_l558 = (! FetchL1Plugin_logic_invalidate_done);
  assign LsuPlugin_logic_frontend_defaultsDecodings_0 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_1 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_2 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_3 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_4 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_5 = 1'b0;
  assign GSharePlugin_logic_mem_writes_0_valid = (GSharePlugin_logic_mem_write_valid && 1'b1);
  assign GSharePlugin_logic_mem_writes_0_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign GSharePlugin_logic_mem_writes_0_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign GSharePlugin_logic_mem_writes_0_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign GSharePlugin_logic_mem_writes_0_payload_data_2 = GSharePlugin_logic_mem_write_payload_data_2;
  assign GSharePlugin_logic_mem_writes_0_payload_data_3 = GSharePlugin_logic_mem_write_payload_data_3;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_0_down_Fetch_WORD_PC[4 : 3];
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = ({_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[0],_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[1]} ^ _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1);
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2 = GSharePlugin_logic_mem_write_payload_data_2;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3 = GSharePlugin_logic_mem_write_payload_data_3;
  assign _zz_GSharePlugin_logic_readRsp_readed_0_0 = fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  assign _zz_GSharePlugin_logic_readRsp_readed_0_0_1 = GSharePlugin_logic_mem_banks_0_spinal_port1;
  assign GSharePlugin_logic_readRsp_readed_0_0 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[1 : 0];
  assign GSharePlugin_logic_readRsp_readed_0_1 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[3 : 2];
  assign GSharePlugin_logic_readRsp_readed_0_2 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[5 : 4];
  assign GSharePlugin_logic_readRsp_readed_0_3 = _zz_GSharePlugin_logic_readRsp_readed_0_0_1[7 : 6];
  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = GSharePlugin_logic_readRsp_readed_0_0;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = GSharePlugin_logic_readRsp_readed_0_1;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 = GSharePlugin_logic_readRsp_readed_0_2;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 = GSharePlugin_logic_readRsp_readed_0_3;
    if(when_GSharePlugin_l100) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3;
    end
  end

  assign when_GSharePlugin_l100 = (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid && (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address == fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH));
  always @(*) begin
    BtbPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(BtbPlugin_logic_applyIt_rasLogic_pushValid) begin
      BtbPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_BtbPlugin_l246) begin
      BtbPlugin_logic_ras_ptr_popIt = 1'b1;
    end
  end

  assign BtbPlugin_logic_ras_write_valid = BtbPlugin_logic_ras_ptr_pushIt;
  assign BtbPlugin_logic_ras_write_payload_address = BtbPlugin_logic_ras_ptr_push;
  always @(*) begin
    BtbPlugin_logic_ras_write_payload_data = 31'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    BtbPlugin_logic_ras_write_payload_data = (_zz_BtbPlugin_logic_ras_write_payload_data >>> 1'd1);
  end

  assign BtbPlugin_logic_memDp_wp_valid = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_memDp_wp_payload_address = BtbPlugin_logic_memWrite_payload_address;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_hash = BtbPlugin_logic_memWrite_payload_data_0_hash;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_sliceLow = BtbPlugin_logic_memWrite_payload_data_0_sliceLow;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget = BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isBranch = BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPush = BtbPlugin_logic_memWrite_payload_data_0_isPush;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPop = BtbPlugin_logic_memWrite_payload_data_0_isPop;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_hash = BtbPlugin_logic_memWrite_payload_data_1_hash;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_sliceLow = BtbPlugin_logic_memWrite_payload_data_1_sliceLow;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_pcTarget = BtbPlugin_logic_memWrite_payload_data_1_pcTarget;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_isBranch = BtbPlugin_logic_memWrite_payload_data_1_isBranch;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_isPush = BtbPlugin_logic_memWrite_payload_data_1_isPush;
  assign BtbPlugin_logic_memDp_wp_payload_data_1_isPop = BtbPlugin_logic_memWrite_payload_data_1_isPop;
  assign BtbPlugin_logic_memDp_wp_payload_mask = BtbPlugin_logic_memWrite_payload_mask;
  assign _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash = BtbPlugin_logic_mem_spinal_port1;
  assign _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1 = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[46 : 0];
  assign _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[93 : 47];
  assign BtbPlugin_logic_memDp_rp_rsp_0_hash = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[11 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_0_sliceLow = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[12 : 12];
  assign BtbPlugin_logic_memDp_rp_rsp_0_pcTarget = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[43 : 13];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isBranch = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[44];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPush = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[45];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPop = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash_1[46];
  assign BtbPlugin_logic_memDp_rp_rsp_1_hash = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[11 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_1_sliceLow = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[12 : 12];
  assign BtbPlugin_logic_memDp_rp_rsp_1_pcTarget = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[43 : 13];
  assign BtbPlugin_logic_memDp_rp_rsp_1_isBranch = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[44];
  assign BtbPlugin_logic_memDp_rp_rsp_1_isPush = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[45];
  assign BtbPlugin_logic_memDp_rp_rsp_1_isPop = _zz_BtbPlugin_logic_memDp_rp_rsp_1_hash[46];
  assign BtbPlugin_logic_memDp_rp_cmd_valid = BtbPlugin_logic_memRead_cmd_valid;
  assign BtbPlugin_logic_memDp_rp_cmd_payload = BtbPlugin_logic_memRead_cmd_payload;
  assign BtbPlugin_logic_memRead_rsp_0_hash = BtbPlugin_logic_memDp_rp_rsp_0_hash;
  assign BtbPlugin_logic_memRead_rsp_0_sliceLow = BtbPlugin_logic_memDp_rp_rsp_0_sliceLow;
  assign BtbPlugin_logic_memRead_rsp_0_pcTarget = BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  assign BtbPlugin_logic_memRead_rsp_0_isBranch = BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  assign BtbPlugin_logic_memRead_rsp_0_isPush = BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  assign BtbPlugin_logic_memRead_rsp_0_isPop = BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  assign BtbPlugin_logic_memRead_rsp_1_hash = BtbPlugin_logic_memDp_rp_rsp_1_hash;
  assign BtbPlugin_logic_memRead_rsp_1_sliceLow = BtbPlugin_logic_memDp_rp_rsp_1_sliceLow;
  assign BtbPlugin_logic_memRead_rsp_1_pcTarget = BtbPlugin_logic_memDp_rp_rsp_1_pcTarget;
  assign BtbPlugin_logic_memRead_rsp_1_isBranch = BtbPlugin_logic_memDp_rp_rsp_1_isBranch;
  assign BtbPlugin_logic_memRead_rsp_1_isPush = BtbPlugin_logic_memDp_rp_rsp_1_isPush;
  assign BtbPlugin_logic_memRead_rsp_1_isPop = BtbPlugin_logic_memDp_rp_rsp_1_isPop;
  assign WhiteboxerPlugin_logic_fetch_fetchId = fetch_logic_ctrls_0_down_Fetch_ID;
  assign WhiteboxerPlugin_logic_decodes_0_fire = ((decode_ctrls_0_up_LANE_SEL_0 && decode_ctrls_0_up_isReady) && (! decode_ctrls_0_lane0_upIsCancel));
  assign when_CtrlLaneApi_l50 = (decode_ctrls_0_up_isReady || decode_ctrls_0_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_0_spawn = (decode_ctrls_0_up_LANE_SEL_0 && (! decode_ctrls_0_up_LANE_SEL_0_regNext));
  assign WhiteboxerPlugin_logic_decodes_0_pc = _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  assign WhiteboxerPlugin_logic_decodes_0_fetchId = decode_ctrls_0_down_Fetch_ID_0;
  assign WhiteboxerPlugin_logic_decodes_0_decodeId = decode_ctrls_0_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_decodes_1_fire = ((decode_ctrls_0_up_LANE_SEL_1 && decode_ctrls_0_up_isReady) && (! decode_ctrls_0_lane1_upIsCancel));
  assign when_CtrlLaneApi_l50_1 = (decode_ctrls_0_up_isReady || decode_ctrls_0_lane1_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_1_spawn = (decode_ctrls_0_up_LANE_SEL_1 && (! decode_ctrls_0_up_LANE_SEL_1_regNext));
  assign WhiteboxerPlugin_logic_decodes_1_pc = _zz_WhiteboxerPlugin_logic_decodes_1_pc;
  assign WhiteboxerPlugin_logic_decodes_1_fetchId = decode_ctrls_0_down_Fetch_ID_1;
  assign WhiteboxerPlugin_logic_decodes_1_decodeId = decode_ctrls_0_down_Decode_DOP_ID_1;
  always @(*) begin
    early0_EnvPlugin_logic_flushPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_flushPort_valid = 1'b1;
    end
  end

  assign early0_EnvPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_trapPort_valid = 1'b1;
    end
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_exception = 1'b1;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_trapPort_payload_tval = ((execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_EBREAK) ? execute_ctrl2_down_PC_lane0 : 32'h0);
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0011;
      end
      EnvPluginOp_ECALL : begin
        early0_EnvPlugin_logic_trapPort_payload_code = (_zz_early0_EnvPlugin_logic_trapPort_payload_code | 4'b1000);
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0001;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b1000;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_arg = 2'bxx;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_arg[1 : 0] = early0_EnvPlugin_logic_exe_xretPriv;
        end
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_trapPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = CsrAccessPlugin_bus_decode_address[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (CsrAccessPlugin_bus_decode_address[11 : 10] == 2'b11);
  assign when_PrivilegedPlugin_l701 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && CsrAccessPlugin_bus_decode_write) || (PrivilegedPlugin_logic_harts_0_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  assign FetchL1Plugin_pmaBuilder_addressBits = FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit[0];
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit = (|1'b1);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_hit = (FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit && FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit);
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = ((FetchL1Plugin_pmaBuilder_addressBits & 32'h80000000) == 32'h80000000);
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = (! ((|{_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault,((FetchL1Plugin_pmaBuilder_addressBits & 32'hf0000000) == 32'h10000000)}) && (|FetchL1Plugin_pmaBuilder_onTransfers_0_hit)));
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = (! _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io[0]);
  assign FetchL1Plugin_logic_bus_toWishbone_pending = (FetchL1Plugin_logic_bus_toWishbone_counter != 1'b0);
  assign FetchL1Plugin_logic_bus_toWishbone_lastCycle = (&FetchL1Plugin_logic_bus_toWishbone_counter);
  assign FetchL1WishbonePlugin_logic_bus_ADR = {_zz_FetchL1WishbonePlugin_logic_bus_ADR,FetchL1Plugin_logic_bus_toWishbone_counter};
  assign FetchL1WishbonePlugin_logic_bus_CTI = (FetchL1Plugin_logic_bus_toWishbone_lastCycle ? 3'b111 : 3'b010);
  assign FetchL1WishbonePlugin_logic_bus_BTE = 2'b00;
  assign FetchL1WishbonePlugin_logic_bus_SEL = 32'hffffffff;
  assign FetchL1WishbonePlugin_logic_bus_WE = 1'b0;
  assign FetchL1WishbonePlugin_logic_bus_DAT_MOSI = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  always @(*) begin
    FetchL1WishbonePlugin_logic_bus_CYC = 1'b0;
    if(when_FetchL1Bus_l247) begin
      FetchL1WishbonePlugin_logic_bus_CYC = 1'b1;
    end
  end

  always @(*) begin
    FetchL1WishbonePlugin_logic_bus_STB = 1'b0;
    if(when_FetchL1Bus_l247) begin
      FetchL1WishbonePlugin_logic_bus_STB = 1'b1;
    end
  end

  assign when_FetchL1Bus_l247 = (FetchL1Plugin_logic_bus_cmd_valid || FetchL1Plugin_logic_bus_toWishbone_pending);
  assign when_FetchL1Bus_l250 = (FetchL1WishbonePlugin_logic_bus_ACK || FetchL1WishbonePlugin_logic_bus_ERR);
  assign FetchL1Plugin_logic_bus_cmd_ready = ((FetchL1Plugin_logic_bus_cmd_valid && FetchL1Plugin_logic_bus_toWishbone_lastCycle) && (FetchL1WishbonePlugin_logic_bus_ACK || FetchL1WishbonePlugin_logic_bus_ERR));
  assign FetchL1Plugin_logic_bus_rsp_valid = _zz_FetchL1Plugin_logic_bus_rsp_valid;
  assign FetchL1Plugin_logic_bus_rsp_payload_id = FetchL1Plugin_logic_bus_cmd_payload_id_regNext;
  assign FetchL1Plugin_logic_bus_rsp_payload_data = FetchL1WishbonePlugin_logic_bus_DAT_MISO_regNext;
  assign FetchL1Plugin_logic_bus_rsp_payload_error = FetchL1WishbonePlugin_logic_bus_ERR_regNext;
  always @(*) begin
    DecoderPlugin_logic_forgetPort_valid = 1'b0;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (decode_ctrls_1_down_PC_0 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice);
    end
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (decode_ctrls_1_down_PC_1 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3);
    end
  end

  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl1_down_integer_RS1_lane0;
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 12],12'h0};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_PC_lane0;
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    early0_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
    if(execute_ctrl2_down_SrcStageables_REVERT_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
    end
    if(execute_ctrl2_down_SrcStageables_ZERO_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1));
  assign execute_ctrl2_down_early0_SrcPlugin_LESS_lane0 = ((execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31] == execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31]) ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0[31] : (execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 ? execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31] : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]));
  assign lane0_IntFormatPlugin_logic_stages_0_hits = {early0_BarrelShifterPlugin_logic_wb_valid,early0_IntAluPlugin_logic_wb_valid};
  assign lane0_IntFormatPlugin_logic_stages_0_wb_valid = (execute_ctrl2_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_0_hits));
  assign lane0_IntFormatPlugin_logic_stages_0_raw = ((lane0_IntFormatPlugin_logic_stages_0_hits[0] ? early0_IntAluPlugin_logic_wb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_0_hits[1] ? early0_BarrelShifterPlugin_logic_wb_payload : 32'h0));
  assign lane0_IntFormatPlugin_logic_stages_0_wb_payload = lane0_IntFormatPlugin_logic_stages_0_raw;
  assign lane0_IntFormatPlugin_logic_stages_1_hits = {LsuPlugin_logic_iwb_valid,{FpuF2iPlugin_logic_iwb_valid,{late0_BarrelShifterPlugin_logic_wb_valid,{late0_IntAluPlugin_logic_wb_valid,early0_MulPlugin_logic_formatBus_valid}}}};
  assign lane0_IntFormatPlugin_logic_stages_1_wb_valid = (execute_ctrl4_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_1_hits));
  assign lane0_IntFormatPlugin_logic_stages_1_raw = ((((lane0_IntFormatPlugin_logic_stages_1_hits[0] ? early0_MulPlugin_logic_formatBus_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_1_hits[1] ? late0_IntAluPlugin_logic_wb_payload : 32'h0)) | ((lane0_IntFormatPlugin_logic_stages_1_hits[2] ? late0_BarrelShifterPlugin_logic_wb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_1_hits[3] ? FpuF2iPlugin_logic_iwb_payload : 32'h0))) | (lane0_IntFormatPlugin_logic_stages_1_hits[4] ? LsuPlugin_logic_iwb_payload : 32'h0));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_1_wb_payload = lane0_IntFormatPlugin_logic_stages_1_raw;
    if(lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[15 : 8] = {8{lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value}};
    end
    if(lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[31 : 16] = {16{lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b01);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1 = lane0_IntFormatPlugin_logic_stages_1_raw[15];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
      end
      2'b01 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b10);
  assign lane0_IntFormatPlugin_logic_stages_2_hits = {FpuMvPlugin_logic_iwb_valid,{FpuCmpPlugin_logic_iwb_valid,{FpuClassPlugin_logic_iwb_valid,{CsrAccessPlugin_logic_wbWi_valid,early0_DivPlugin_logic_formatBus_valid}}}};
  assign lane0_IntFormatPlugin_logic_stages_2_wb_valid = (execute_ctrl3_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_2_hits));
  assign lane0_IntFormatPlugin_logic_stages_2_raw = ((((lane0_IntFormatPlugin_logic_stages_2_hits[0] ? early0_DivPlugin_logic_formatBus_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[1] ? CsrAccessPlugin_logic_wbWi_payload : 32'h0)) | ((lane0_IntFormatPlugin_logic_stages_2_hits[2] ? FpuClassPlugin_logic_iwb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[3] ? FpuCmpPlugin_logic_iwb_payload : 32'h0))) | (lane0_IntFormatPlugin_logic_stages_2_hits[4] ? FpuMvPlugin_logic_iwb_payload : 32'h0));
  assign lane0_IntFormatPlugin_logic_stages_2_wb_payload = lane0_IntFormatPlugin_logic_stages_2_raw;
  always @(*) begin
    _zz_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = execute_ctrl3_down_integer_RS1_lane0;
      end
      default : begin
        _zz_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = {execute_ctrl3_down_Decode_UOP_lane0[31 : 12],12'h0};
      end
    endcase
  end

  assign execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = _zz_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = execute_ctrl3_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = execute_ctrl3_down_PC_lane0;
      end
      default : begin
      end
    endcase
  end

  assign execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = _zz_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    late0_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0;
    if(execute_ctrl4_down_SrcStageables_REVERT_lane0) begin
      late0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
    end
    if(execute_ctrl4_down_SrcStageables_ZERO_lane0) begin
      late0_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1));
  assign execute_ctrl4_down_late0_SrcPlugin_LESS_lane0 = ((execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31] == execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[31]) ? execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0[31] : (execute_ctrl4_down_SrcStageables_UNSIGNED_lane0 ? execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[31] : execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]));
  always @(*) begin
    _zz_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1)
      1'b0 : begin
        _zz_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = execute_ctrl1_down_integer_RS1_lane1;
      end
      default : begin
        _zz_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = {execute_ctrl1_down_Decode_UOP_lane1[31 : 12],12'h0};
      end
    endcase
  end

  assign execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = _zz_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  always @(*) begin
    _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1)
      2'b00 : begin
        _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = execute_ctrl1_down_integer_RS2_lane1;
      end
      2'b01 : begin
        _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = {{20{_zz__zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1[11]}}, _zz__zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1};
      end
      2'b10 : begin
        _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = execute_ctrl1_down_PC_lane1;
      end
      default : begin
      end
    endcase
  end

  assign execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = _zz_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  always @(*) begin
    early1_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1;
    if(execute_ctrl2_down_SrcStageables_REVERT_lane1) begin
      early1_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
    end
    if(execute_ctrl2_down_SrcStageables_ZERO_lane1) begin
      early1_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 = ($signed(_zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1) + $signed(_zz_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1));
  assign execute_ctrl2_down_early1_SrcPlugin_LESS_lane1 = ((execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31] == execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[31]) ? execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1[31] : (execute_ctrl2_down_SrcStageables_UNSIGNED_lane1 ? execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[31] : execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]));
  assign lane1_IntFormatPlugin_logic_stages_0_hits = {early1_BarrelShifterPlugin_logic_wb_valid,early1_IntAluPlugin_logic_wb_valid};
  assign lane1_IntFormatPlugin_logic_stages_0_wb_valid = (execute_ctrl2_up_LANE_SEL_lane1 && (|lane1_IntFormatPlugin_logic_stages_0_hits));
  assign lane1_IntFormatPlugin_logic_stages_0_raw = ((lane1_IntFormatPlugin_logic_stages_0_hits[0] ? early1_IntAluPlugin_logic_wb_payload : 32'h0) | (lane1_IntFormatPlugin_logic_stages_0_hits[1] ? early1_BarrelShifterPlugin_logic_wb_payload : 32'h0));
  assign lane1_IntFormatPlugin_logic_stages_0_wb_payload = lane1_IntFormatPlugin_logic_stages_0_raw;
  assign lane1_IntFormatPlugin_logic_stages_1_hits = {late1_BarrelShifterPlugin_logic_wb_valid,late1_IntAluPlugin_logic_wb_valid};
  assign lane1_IntFormatPlugin_logic_stages_1_wb_valid = (execute_ctrl4_up_LANE_SEL_lane1 && (|lane1_IntFormatPlugin_logic_stages_1_hits));
  assign lane1_IntFormatPlugin_logic_stages_1_raw = ((lane1_IntFormatPlugin_logic_stages_1_hits[0] ? late1_IntAluPlugin_logic_wb_payload : 32'h0) | (lane1_IntFormatPlugin_logic_stages_1_hits[1] ? late1_BarrelShifterPlugin_logic_wb_payload : 32'h0));
  assign lane1_IntFormatPlugin_logic_stages_1_wb_payload = lane1_IntFormatPlugin_logic_stages_1_raw;
  always @(*) begin
    _zz_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1)
      1'b0 : begin
        _zz_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = execute_ctrl3_down_integer_RS1_lane1;
      end
      default : begin
        _zz_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = {execute_ctrl3_down_Decode_UOP_lane1[31 : 12],12'h0};
      end
    endcase
  end

  assign execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = _zz_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  always @(*) begin
    _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1)
      2'b00 : begin
        _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = execute_ctrl3_down_integer_RS2_lane1;
      end
      2'b01 : begin
        _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = {{20{_zz__zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1[11]}}, _zz__zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1};
      end
      2'b10 : begin
        _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = execute_ctrl3_down_PC_lane1;
      end
      default : begin
      end
    endcase
  end

  assign execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = _zz_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  always @(*) begin
    late1_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1;
    if(execute_ctrl4_down_SrcStageables_REVERT_lane1) begin
      late1_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
    end
    if(execute_ctrl4_down_SrcStageables_ZERO_lane1) begin
      late1_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 = ($signed(_zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1) + $signed(_zz_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1));
  assign execute_ctrl4_down_late1_SrcPlugin_LESS_lane1 = ((execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31] == execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[31]) ? execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1[31] : (execute_ctrl4_down_SrcStageables_UNSIGNED_lane1 ? execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[31] : execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]));
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode = FpuAddPlugin_logic_addPort_cmd_rs1_mode;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_0_quiet = FpuAddPlugin_logic_addPort_cmd_rs1_quiet;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_0_sign = FpuAddPlugin_logic_addPort_cmd_rs1_sign;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent = _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_0_mantissa = ({53'd0,FpuAddPlugin_logic_addPort_cmd_rs1_mantissa} <<< 6'd53);
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode = FpuMulPlugin_logic_addPort_cmd_rs1_mode;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_1_quiet = FpuMulPlugin_logic_addPort_cmd_rs1_quiet;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_1_sign = FpuMulPlugin_logic_addPort_cmd_rs1_sign;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent = _zz_FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent;
  assign FpuAddSharedPlugin_logic_inserter_portsRs1_1_mantissa = FpuMulPlugin_logic_addPort_cmd_rs1_mantissa;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode = FpuAddPlugin_logic_addPort_cmd_rs2_mode;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_0_quiet = FpuAddPlugin_logic_addPort_cmd_rs2_quiet;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_0_sign = FpuAddPlugin_logic_addPort_cmd_rs2_sign;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent = _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_0_mantissa = FpuAddPlugin_logic_addPort_cmd_rs2_mantissa;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode = FpuMulPlugin_logic_addPort_cmd_rs2_mode;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_1_quiet = FpuMulPlugin_logic_addPort_cmd_rs2_quiet;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_1_sign = FpuMulPlugin_logic_addPort_cmd_rs2_sign;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent = _zz_FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent;
  assign FpuAddSharedPlugin_logic_inserter_portsRs2_1_mantissa = FpuMulPlugin_logic_addPort_cmd_rs2_mantissa;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_valid = (|FpuAddPlugin_logic_addPort_cmd_at);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1 = (|FpuMulPlugin_logic_addPort_cmd_at);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet = {_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1,_zz_FpuAddSharedPlugin_logic_pip_node_0_valid};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1 = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet[0] ? {FpuAddSharedPlugin_logic_inserter_portsRs1_0_mantissa,{FpuAddSharedPlugin_logic_inserter_portsRs1_0_exponent,{FpuAddSharedPlugin_logic_inserter_portsRs1_0_sign,{FpuAddSharedPlugin_logic_inserter_portsRs1_0_quiet,FpuAddSharedPlugin_logic_inserter_portsRs1_0_mode}}}} : 122'h0) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet[1] ? {FpuAddSharedPlugin_logic_inserter_portsRs1_1_mantissa,{FpuAddSharedPlugin_logic_inserter_portsRs1_1_exponent,{FpuAddSharedPlugin_logic_inserter_portsRs1_1_sign,{FpuAddSharedPlugin_logic_inserter_portsRs1_1_quiet,FpuAddSharedPlugin_logic_inserter_portsRs1_1_mode}}}} : 122'h0));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1 = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1[1 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode_1;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1[2];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_sign = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet_1[3];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_exponent;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa[104 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet = {_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1,_zz_FpuAddSharedPlugin_logic_pip_node_0_valid};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1 = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet[0] ? {FpuAddSharedPlugin_logic_inserter_portsRs2_0_mantissa,{FpuAddSharedPlugin_logic_inserter_portsRs2_0_exponent,{FpuAddSharedPlugin_logic_inserter_portsRs2_0_sign,{FpuAddSharedPlugin_logic_inserter_portsRs2_0_quiet,FpuAddSharedPlugin_logic_inserter_portsRs2_0_mode}}}} : 68'h0) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet[1] ? {FpuAddSharedPlugin_logic_inserter_portsRs2_1_mantissa,{FpuAddSharedPlugin_logic_inserter_portsRs2_1_exponent,{FpuAddSharedPlugin_logic_inserter_portsRs2_1_sign,{FpuAddSharedPlugin_logic_inserter_portsRs2_1_quiet,FpuAddSharedPlugin_logic_inserter_portsRs2_1_mode}}}} : 68'h0));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1 = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1[1 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode_1;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1[2];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_sign = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet_1[3];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_exponent;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa[51 : 0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1 = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_valid ? FpuAddPlugin_logic_addPort_cmd_format : 1'b0) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1 ? FpuMulPlugin_logic_addPort_cmd_format : 1'b0));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT_1;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1 = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_valid ? FpuAddPlugin_logic_addPort_cmd_roundMode : 3'b000) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1 ? FpuMulPlugin_logic_addPort_cmd_roundMode : 3'b000));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE_1;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE;
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_RDN = (FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE == FpuRoundMode_RDN);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_valid ? {FpuAddPlugin_logic_addPort_cmd_flags_NV,{FpuAddPlugin_logic_addPort_cmd_flags_DZ,{FpuAddPlugin_logic_addPort_cmd_flags_OF,{FpuAddPlugin_logic_addPort_cmd_flags_UF,FpuAddPlugin_logic_addPort_cmd_flags_NX}}}} : 5'h0) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1 ? {FpuMulPlugin_logic_addPort_cmd_flags_NV,{FpuMulPlugin_logic_addPort_cmd_flags_DZ,{FpuMulPlugin_logic_addPort_cmd_flags_OF,{FpuMulPlugin_logic_addPort_cmd_flags_UF,FpuMulPlugin_logic_addPort_cmd_flags_NX}}}} : 5'h0));
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX[0];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_UF = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX[1];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_OF = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX[2];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_DZ = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX[3];
  assign FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NV = _zz_FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX[4];
  assign FpuAddSharedPlugin_logic_pip_node_0_Decode_UOP_ID = ((_zz_FpuAddSharedPlugin_logic_pip_node_0_valid ? FpuAddPlugin_logic_addPort_cmd_uopId : 16'h0) | (_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1 ? FpuMulPlugin_logic_addPort_cmd_uopId : 16'h0));
  assign FpuAddSharedPlugin_logic_pip_node_0_valid = (|{_zz_FpuAddSharedPlugin_logic_pip_node_0_valid_1,_zz_FpuAddSharedPlugin_logic_pip_node_0_valid});
  always @(*) begin
    FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH[0] = (|FpuAddPlugin_logic_addPort_cmd_at[0]);
    FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH[1] = (|FpuMulPlugin_logic_addPort_cmd_at[0]);
  end

  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21 = _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21;
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12 = _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp12;
  assign _zz_when_AFix_l1168 = (FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21[12] ? _zz__zz_when_AFix_l1168 : _zz__zz_when_AFix_l1168_1);
  assign when_AFix_l1168 = _zz_when_AFix_l1168[12];
  always @(*) begin
    if(when_AFix_l1168) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs = 13'h0;
    end else begin
      _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs = _zz_when_AFix_l1168;
    end
  end

  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs = _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs[11 : 0];
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentBigger = ((FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_exp21[12] || (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode == FloatMode_ZERO)) && (! (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode == FloatMode_ZERO)));
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual = ($signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual) == $signed(_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual_1));
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger = (_zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger < FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa);
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_absRs1Bigger = ((((FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentBigger || (FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1ExponentEqual && FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_rs1MantissaBigger)) && (! (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode == FloatMode_ZERO))) || (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode == FloatMode_INF)) && (! (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode == FloatMode_INF)));
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_needSub = (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_sign ^ FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_sign);
  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_passThrough = ((FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode == FloatMode_ZERO) || (FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode == FloatMode_ZERO));
  assign when_UInt_l119 = (|FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs[11 : 7]);
  always @(*) begin
    if(when_UInt_l119) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat = 7'h7f;
    end else begin
      _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat = FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbs[6 : 0];
    end
  end

  assign FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat = (FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_passThrough ? 7'h7f : _zz_FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat);
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xySign = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger ? FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_sign : FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_sign);
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa = _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa;
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted = _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted;
  assign _zz_when_Utils_l1585_14 = {{FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissaUnshifted,1'b0},1'b0};
  always @(*) begin
    _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b0;
    if(when_Utils_l1585) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_1) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_2) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_3) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_4) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_5) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
    if(when_Utils_l1585_6) begin
      _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_1 = 1'b1;
    end
  end

  assign when_Utils_l1585 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[0] && (_zz_when_Utils_l1585_14[0 : 0] != 1'b0));
  assign when_Utils_l1585_1 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[1] && (_zz_when_Utils_l1585_13[1 : 0] != 2'b00));
  assign when_Utils_l1585_2 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[2] && (_zz_when_Utils_l1585_12[3 : 0] != 4'b0000));
  assign when_Utils_l1585_3 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[3] && (_zz_when_Utils_l1585_11[7 : 0] != 8'h0));
  assign when_Utils_l1585_4 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[4] && (_zz_when_Utils_l1585_10[15 : 0] != 16'h0));
  assign when_Utils_l1585_5 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[5] && (_zz_when_Utils_l1585_9[31 : 0] != 32'h0));
  assign when_Utils_l1585_6 = (FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat[6] && (_zz_when_Utils_l1585_8[63 : 0] != 64'h0));
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter = (_zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter | _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter_2);
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissa = FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter[107 : 1];
  assign FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent = _zz_FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xyExponent;
  always @(*) begin
    FpuAddSharedPlugin_logic_pip_node_2_adder_math_roundingScrap = (FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_shifter[0] && (! FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_passThrough));
    if(when_FpuAdd_l56) begin
      FpuAddSharedPlugin_logic_pip_node_2_adder_math_roundingScrap = 1'b0;
    end
  end

  assign when_FpuAdd_l56 = ((! (FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode == FloatMode_NORMAL)) || (! (FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode == FloatMode_NORMAL)));
  assign _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned = FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_yMantissa;
  assign FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned = _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_ySigned_1;
  assign FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa = _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa[107:0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh = {FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[0],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[1],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[2],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[3],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[4],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[5],{FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa[6],{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh,{_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1,_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2}}}}}}}}};
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[0];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[1];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[2];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[3];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[4];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[5];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[6];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[7];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[8];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[9];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[10];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[11];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[12];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[13];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[14];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[15];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[16];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[17];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[18];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[19];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[20];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[21];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[22];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[23];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[24];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[25];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[26];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[27];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[28];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[29];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_31 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[30];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_32 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[31];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[32];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[33];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_35 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[34];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_36 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[35];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[36];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[37];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_39 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[38];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_40 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[39];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[40];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[41];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_43 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[42];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_44 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[43];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[44];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[45];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_47 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[46];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_48 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[47];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[48];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[49];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_51 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[50];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_52 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[51];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[52];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[53];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_55 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[54];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_56 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[55];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[56];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[57];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_59 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[58];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_60 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[59];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[60];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[61];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_63 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[62];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_64 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[63];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[64];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[65];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_67 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[66];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_68 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[67];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[68];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[69];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_71 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[70];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_72 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[71];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[72];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[73];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_75 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[74];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_76 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[75];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[76];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[77];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_79 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[78];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_80 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[79];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[80];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[81];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_83 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[82];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_84 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[83];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[84];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[85];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_87 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[86];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_88 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[87];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[88];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[89];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_91 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[90];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_92 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[91];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[92];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[93];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_95 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[94];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_96 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[95];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[96];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[97];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_99 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[98];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_100 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[99];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[100];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[101];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_103 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[102];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_104 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[103];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[104];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_106 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[105];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_107 = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[106];
  always @(*) begin
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[0] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1 && (! 1'b0));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[1] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2 && (! _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[2] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3 && (! (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1})));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[3] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4 && (! (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1}})));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[4] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5 && (! _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[5] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[6] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[7] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5}}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[8] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[9] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[10] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[11] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9}}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[12] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_112 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[13] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[14] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[15] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13}}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[16] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_114 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[17] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[18] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[19] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17}}) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[20] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115)));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[21] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[22] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[23] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[24] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[25] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[26] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[27] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[28] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_119 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[29] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[30] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_31 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[31] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_32 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_31,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[32] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_121 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[33] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[34] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_35 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[35] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_36 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_35,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[36] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[37] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[38] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_39 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[39] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_40 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_39,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[40] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[41] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[42] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_43 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[43] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_44 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_43,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[44] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_127 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[45] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[46] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_47 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[47] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_48 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_47,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[48] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_129 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[49] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[50] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_51 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[51] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_52 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_51,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[52] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[53] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[54] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_55 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[55] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_56 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_55,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[56] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[57] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[58] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_59 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[59] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_60 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_59,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[60] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_135 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[61] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[62] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_63 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[63] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_64 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_63,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[64] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_137 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[65] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[66] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_67 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[67] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_68 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_67,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[68] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[69] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[70] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_71 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[71] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_72 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_71,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[72] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[73] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[74] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_75 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[75] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_76 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_75,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[76] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_143 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[77] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[78] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_79 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[79] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_80 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_79,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[80] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_145 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[81] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[82] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_83 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[83] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_84 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_83,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[84] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[85] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[86] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_87 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[87] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_88 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_87,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[88] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[89] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[90] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_91 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[91] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_92 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_91,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[92] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_150 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[93] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[94] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_95 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[95] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_96 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_95,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[96] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_152 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[97] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[98] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_99 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[99] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_100 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_99,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[100] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[101] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[102] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_103 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[103] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_104 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_103,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[104] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_156 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[105] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_106 && (! (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_157 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[106] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_107 && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_106,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_157 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
    _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108[107] = (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[107] && (! ((|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_107,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_106,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_105}}) || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_157 || (_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140)))));
  end

  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_4,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_3,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_2,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_1}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_8,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_7,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_6,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_5}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_111 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_112 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_12,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_11,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_10,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_9}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_113 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_112,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_114 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_16,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_15,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_14,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_13}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_114,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_112,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_110,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_109}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_20,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_19,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_18,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_17}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_24,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_23,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_22,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_21}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_118 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_119 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_28,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_27,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_26,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_25}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_120 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_119,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_121 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_32,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_31,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_30,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_29}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_121,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_119,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_117,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_116}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_36,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_35,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_34,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_33}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_124 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_40,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_39,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_38,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_37}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_126 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_127 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_44,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_43,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_42,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_41}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_128 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_127,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_129 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_48,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_47,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_46,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_45}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_129,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_127,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_125,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_123}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_52,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_51,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_50,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_49}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_132 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_56,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_55,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_54,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_53}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_134 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_135 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_60,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_59,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_58,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_57}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_136 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_135,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_137 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_64,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_63,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_62,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_61}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_137,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_135,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_133,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_131}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_68,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_67,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_66,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_65}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_140 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_138,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_130,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_122,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_115}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_72,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_71,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_70,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_69}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_142 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_143 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_76,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_75,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_74,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_73}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_144 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_143,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_145 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_80,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_79,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_78,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_77}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_145,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_143,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_141,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_139}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_84,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_83,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_82,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_81}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_88,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_87,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_86,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_85}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_149 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_150 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_92,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_91,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_90,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_89}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_151 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_150,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_152 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_96,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_95,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_94,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_93}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_152,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_150,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_148,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_147}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_100,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_99,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_98,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_97}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_155 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_153,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_146});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_156 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_104,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_103,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_102,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_101}}});
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_157 = (|{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_156,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_154});
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh = _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh_108;
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[3];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_1 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[5];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_2 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[6];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_3 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[7];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_4 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[9];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_5 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[10];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_6 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[11];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_7 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[12];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_8 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[13];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_9 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[14];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_10 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[15];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_11 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[17];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_12 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[18];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_13 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[19];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_14 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[20];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_15 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[21];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_16 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[22];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_17 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[23];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_18 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[24];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_19 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[25];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_20 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[26];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_21 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[27];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_22 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[28];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_23 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[29];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_24 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[30];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_25 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[31];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_26 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[33];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_27 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[34];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_28 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[35];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_29 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[36];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_30 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[37];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_31 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[38];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_32 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[39];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_33 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[40];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_34 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[41];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_35 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[42];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_36 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[43];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_37 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[44];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_38 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[45];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_39 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[46];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_40 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[47];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_41 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[48];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_42 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[49];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_43 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[50];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_44 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[51];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_45 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[52];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_46 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[53];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_47 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[54];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_48 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[55];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_49 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[56];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_50 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[57];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_51 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[58];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_52 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[59];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[60];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[61];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[62];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[63];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_57 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[65];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_58 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[66];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_59 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[67];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_60 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[68];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_61 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[69];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_62 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[70];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[71];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_64 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[72];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_65 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[73];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_66 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[74];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[75];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_68 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[76];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[77];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[78];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[79];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_72 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[80];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_73 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[81];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_74 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[82];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[83];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_76 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[84];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[85];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[86];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[87];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_80 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[88];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[89];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[90];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[91];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[92];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[93];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[94];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[95];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_88 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[96];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_89 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[97];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_90 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[98];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[99];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_92 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[100];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[101];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[102];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[103];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_96 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[104];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[105];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[106];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99 = FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shiftOh[107];
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_73) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_89) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_74) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_90) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_63) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_68) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_76) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_92) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103 = (((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_67) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_68) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_69) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_70) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_71) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_80) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_96) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_72) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_73) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_74) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_75) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_76) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_77) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_78) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_79) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_80) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_81) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_82) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_83) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_53) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_54) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_55) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_56) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_88) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_89) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_90) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_92) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_96) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99);
  assign _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106 = ((((((((((((((((_zz__zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106 || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_84) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_85) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_86) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_87) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_88) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_89) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_90) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_91) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_92) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_93) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_94) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_95) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_96) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_97) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_98) || _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_99);
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift = {_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_106,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_105,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_104,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_103,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_102,{_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_101,_zz_FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift_100}}}}}};
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceInfinity = ((FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode == FloatMode_INF) || (FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode == FloatMode_INF));
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceZero = ((FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa == 108'h0) || ((FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode == FloatMode_ZERO) && (FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode == FloatMode_ZERO)));
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_infinityNan = (((FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode == FloatMode_INF) && (FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode == FloatMode_INF)) && (FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_sign ^ FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_sign));
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceNan = (((FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode == FloatMode_NAN) || (FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode == FloatMode_NAN)) || FpuAddSharedPlugin_logic_pip_node_3_adder_norm_infinityNan);
  assign FpuAddSharedPlugin_logic_pip_node_3_adder_norm_xyMantissaZero = (FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa == 108'h0);
  assign FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_exponent;
  assign FpuAddSharedPlugin_logic_pip_node_4_adder_result_mantissa = (FpuAddSharedPlugin_logic_pip_node_4_adder_math_xyMantissa <<< FpuAddSharedPlugin_logic_pip_node_4_adder_norm_shift);
  always @(*) begin
    FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_sign = FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xySign;
    if(!FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceNan) begin
      if(!FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceInfinity) begin
        if(FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceZero) begin
          if(when_FpuAdd_l101) begin
            FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_sign = (FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_sign && FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_sign);
          end
          if(when_FpuAdd_l104) begin
            FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_sign = 1'b1;
          end
        end
      end
    end
  end

  assign FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa[107:0];
  assign FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent = _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_exponent;
  always @(*) begin
    FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_quiet = 1'b0;
    if(FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceNan) begin
      FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_quiet = 1'b1;
    end
  end

  always @(*) begin
    FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode = FloatMode_NORMAL;
    if(FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceNan) begin
      FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode = FloatMode_NAN;
    end else begin
      if(FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceInfinity) begin
        FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode = FloatMode_INF;
      end else begin
        if(FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceZero) begin
          FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode = FloatMode_ZERO;
        end
      end
    end
  end

  assign FpuAddSharedPlugin_logic_pip_node_4_adder_result_NV = ((FpuAddSharedPlugin_logic_pip_node_4_adder_norm_infinityNan || ((FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode == FloatMode_NAN) && (! FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_quiet))) || ((FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode == FloatMode_NAN) && (! FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_quiet)));
  assign when_FpuAdd_l101 = (FpuAddSharedPlugin_logic_pip_node_4_adder_norm_xyMantissaZero || ((FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode == FloatMode_ZERO) && (FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode == FloatMode_ZERO)));
  assign when_FpuAdd_l104 = ((FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_sign || FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_sign) && FpuAddSharedPlugin_logic_pip_node_4_inserter_RDN);
  assign FpuAddSharedPlugin_logic_onPack_mask = (FpuAddSharedPlugin_logic_pip_node_4_inserter_GROUP_OH & {execute_ctrl9_up_LANE_SEL_lane0,execute_ctrl6_up_LANE_SEL_lane0});
  assign FpuAddSharedPlugin_logic_packPort_cmd_at = FpuAddSharedPlugin_logic_onPack_mask;
  assign FpuAddSharedPlugin_logic_packPort_cmd_value_mode = FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mode;
  assign FpuAddSharedPlugin_logic_packPort_cmd_value_quiet = FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_quiet;
  assign FpuAddSharedPlugin_logic_packPort_cmd_value_sign = FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_sign;
  assign FpuAddSharedPlugin_logic_packPort_cmd_value_exponent = _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_when_AFix_l852 = FpuAddSharedPlugin_logic_pip_node_4_adder_result_RESULT_mantissa;
  always @(*) begin
    _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa = _zz_when_AFix_l852[107 : 54];
    if(when_AFix_l852) begin
      _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa[0] = 1'b1;
    end
  end

  assign when_AFix_l852 = (|_zz_when_AFix_l852[53 : 0]);
  assign FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa = _zz_FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuAddSharedPlugin_logic_packPort_cmd_format = FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT;
  assign FpuAddSharedPlugin_logic_packPort_cmd_roundMode = FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE;
  assign FpuAddSharedPlugin_logic_packPort_cmd_uopId = FpuAddSharedPlugin_logic_pip_node_4_Decode_UOP_ID;
  assign FpuAddSharedPlugin_logic_packPort_cmd_flags_NX = FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NX;
  assign FpuAddSharedPlugin_logic_packPort_cmd_flags_UF = FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_UF;
  assign FpuAddSharedPlugin_logic_packPort_cmd_flags_OF = FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_OF;
  assign FpuAddSharedPlugin_logic_packPort_cmd_flags_DZ = FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_DZ;
  always @(*) begin
    FpuAddSharedPlugin_logic_packPort_cmd_flags_NV = FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NV;
    if(FpuAddSharedPlugin_logic_pip_node_4_adder_result_NV) begin
      FpuAddSharedPlugin_logic_packPort_cmd_flags_NV = 1'b1;
    end
  end

  assign FpuAddSharedPlugin_logic_pip_node_4_ready = (! execute_freeze_valid);
  assign FpuAddSharedPlugin_logic_pip_node_0_ready = FpuAddSharedPlugin_logic_pip_node_1_ready;
  assign FpuAddSharedPlugin_logic_pip_node_1_ready = FpuAddSharedPlugin_logic_pip_node_2_ready;
  assign FpuAddSharedPlugin_logic_pip_node_2_ready = FpuAddSharedPlugin_logic_pip_node_3_ready;
  assign FpuAddSharedPlugin_logic_pip_node_3_ready = FpuAddSharedPlugin_logic_pip_node_4_ready;
  assign FpuAddSharedPlugin_logic_pip_node_0_isValid = FpuAddSharedPlugin_logic_pip_node_0_valid;
  assign FpuAddSharedPlugin_logic_pip_node_0_isReady = FpuAddSharedPlugin_logic_pip_node_0_ready;
  assign FpuAddSharedPlugin_logic_pip_node_1_isValid = FpuAddSharedPlugin_logic_pip_node_1_valid;
  assign FpuAddSharedPlugin_logic_pip_node_1_isReady = FpuAddSharedPlugin_logic_pip_node_1_ready;
  assign FpuAddSharedPlugin_logic_pip_node_2_isValid = FpuAddSharedPlugin_logic_pip_node_2_valid;
  assign FpuAddSharedPlugin_logic_pip_node_2_isReady = FpuAddSharedPlugin_logic_pip_node_2_ready;
  assign FpuAddSharedPlugin_logic_pip_node_3_isValid = FpuAddSharedPlugin_logic_pip_node_3_valid;
  assign FpuAddSharedPlugin_logic_pip_node_3_isReady = FpuAddSharedPlugin_logic_pip_node_3_ready;
  assign FpuUnpackerPlugin_logic_unpacker_node_0_valid = FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_valid;
  assign FpuUnpackerPlugin_logic_unpacker_node_0_input_args_data = FpuUnpackerPlugin_logic_unpacker_arbiter_io_output_payload_data;
  assign FpuUnpackerPlugin_logic_unpacker_node_0_input_source = FpuUnpackerPlugin_logic_unpacker_arbiter_io_chosen;
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy = ({1'd0,{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[0],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[1],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[2],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[3],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[4],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[5],{FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data[6],{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy,{_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1,_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2}}}}}}}}}} <<< 1'd1);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[0];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[1];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[2];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[3];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[4];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[5];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[6];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[7];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[8];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[9];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[10];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_12 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[11];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[12];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[13];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_15 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[14];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_16 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[15];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[16];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[17];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_19 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[18];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_20 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[19];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[20];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[21];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_23 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[22];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_24 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[23];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[24];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[25];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_27 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[26];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_28 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[27];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[28];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[29];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_31 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[30];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_32 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[31];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[32];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[33];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_35 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[34];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_36 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[35];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[36];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[37];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_39 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[38];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_40 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[39];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[40];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[41];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_43 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[42];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_44 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[43];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[44];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[45];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_47 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[46];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_48 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[47];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[48];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[49];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_51 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[50];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_52 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[51];
  always @(*) begin
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[0] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1 && (! 1'b0));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[1] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2 && (! _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[2] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3 && (! (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1})));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[3] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4 && (! (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1}})));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[4] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5 && (! _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[5] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[6] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[7] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5}}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[8] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[9] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[10] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[11] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_12 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9}}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[12] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_57 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[13] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[14] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_15 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[15] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_16 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_15,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13}}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[16] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_59 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[17] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[18] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_19 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[19] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_20 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_19,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17}}) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[20] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60)));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[21] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[22] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_23 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[23] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_24 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_23,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[24] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[25] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[26] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_27 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[27] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_28 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_27,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[28] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_64 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[29] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[30] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_31 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[31] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_32 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_31,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[32] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_66 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[33] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[34] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_35 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[35] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_36 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_35,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[36] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[37] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[38] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_39 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[39] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_40 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_39,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[40] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[41] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[42] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_43 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[43] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_44 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_43,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[44] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_72 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[45] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[46] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_47 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[47] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_48 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_47,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[48] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_74 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[49] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50 && (! (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49 || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[50] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_51 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[51] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_52 && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_51,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
    _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53[52] = (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy[52] && (! ((|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_52,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_51,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_50,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_49}}}) || (_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69))));
  end

  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_4,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_3,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_2,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_1}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_8,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_7,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_6,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_5}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_56 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_57 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_12,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_11,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_10,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_9}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_58 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_57,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_59 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_16,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_15,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_14,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_13}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_59,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_57,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_55,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_54}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_20,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_19,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_18,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_17}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_24,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_23,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_22,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_21}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_63 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_64 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_28,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_27,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_26,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_25}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_65 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_64,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_66 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_32,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_31,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_30,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_29}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_66,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_64,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_62,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_61}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_36,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_35,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_34,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_33}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_69 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_67,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_60});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_40,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_39,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_38,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_37}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_71 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_72 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_44,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_43,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_42,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_41}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_73 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_72,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_74 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_48,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_47,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_46,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_45}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_75 = (|{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_74,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_72,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_70,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_68}}});
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_53;
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_77 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[3];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_78 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[5];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_79 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[6];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_80 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[7];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_81 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[9];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_82 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[10];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_83 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[11];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_84 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[12];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_85 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[13];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_86 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[14];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_87 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[15];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_88 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[17];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_89 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[18];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_90 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[19];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_91 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[20];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_92 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[21];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_93 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[22];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[23];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_95 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[24];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_96 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[25];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_97 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[26];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[27];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_99 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[28];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[29];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[30];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[31];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_103 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[33];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_104 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[34];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_105 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[35];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_106 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[36];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_107 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[37];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_108 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[38];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[39];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_110 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[40];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_111 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[41];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_112 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[42];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[43];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_114 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[44];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[45];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[46];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[47];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_118 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[48];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_119 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[49];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_120 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[50];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[51];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_122 = _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_76[52];
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123 = ((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_92) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_96) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_103) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_105) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_107) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_111) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_119) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124 = ((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_93) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_97) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_104) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_105) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_108) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_112) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_120) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125 = (((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_91) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_92) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_93) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_99) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_106) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_107) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_108) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_114) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_122);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126 = ((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_95) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_96) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_97) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_99) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_110) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_111) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_112) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_114) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127 = ((((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_90) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_91) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_92) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_93) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_94) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_95) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_96) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_97) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_98) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_99) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_100) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_101) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_102) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_118) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_119) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_120) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_122);
  assign _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128 = ((((((((((((((((_zz__zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128 || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_107) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_108) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_109) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_110) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_111) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_112) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_113) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_114) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_115) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_116) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_117) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_118) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_119) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_120) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_121) || _zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_122);
  assign FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy = {_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_128,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_127,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_126,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_125,{_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_124,_zz_FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy_123}}}}};
  assign FpuUnpackerPlugin_logic_unpacker_logic_shifter = (FpuUnpackerPlugin_logic_unpacker_node_2_input_args_data <<< FpuUnpackerPlugin_logic_unpacker_node_2_setup_shiftBy);
  always @(*) begin
    FpuUnpackerPlugin_logic_unpacker_results_0_valid = 1'b0;
    if(FpuUnpackerPlugin_logic_unpacker_node_2_isValid) begin
      if(_zz_46[0]) begin
        FpuUnpackerPlugin_logic_unpacker_results_0_valid = 1'b1;
      end
    end
  end

  assign FpuUnpackerPlugin_logic_unpacker_results_0_payload_data = FpuUnpackerPlugin_logic_unpacker_logic_shifter;
  assign FpuUnpackerPlugin_logic_unpacker_results_0_payload_shift = FpuUnpackerPlugin_logic_unpacker_node_2_setup_shiftBy;
  always @(*) begin
    FpuUnpackerPlugin_logic_unpacker_results_1_valid = 1'b0;
    if(FpuUnpackerPlugin_logic_unpacker_node_2_isValid) begin
      if(_zz_46[1]) begin
        FpuUnpackerPlugin_logic_unpacker_results_1_valid = 1'b1;
      end
    end
  end

  assign FpuUnpackerPlugin_logic_unpacker_results_1_payload_data = FpuUnpackerPlugin_logic_unpacker_logic_shifter;
  assign FpuUnpackerPlugin_logic_unpacker_results_1_payload_shift = FpuUnpackerPlugin_logic_unpacker_node_2_setup_shiftBy;
  assign _zz_46 = ({1'd0,1'b1} <<< FpuUnpackerPlugin_logic_unpacker_node_2_input_source);
  always @(*) begin
    FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid = 1'b0;
    if(when_FpuUnpackerPlugin_l243) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid = 1'b1;
    end
    if(when_FpuUnpackerPlugin_l243_1) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid = 1'b1;
    end
    if(when_FpuUnpackerPlugin_l243_2) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_valid = 1'b1;
    end
  end

  always @(*) begin
    FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_FpuUnpackerPlugin_l243) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa;
    end
    if(when_FpuUnpackerPlugin_l243_1) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa;
    end
    if(when_FpuUnpackerPlugin_l243_2) begin
      FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_0_payload_data = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa;
    end
  end

  assign when_FpuUnpackerPlugin_l165 = (! execute_freeze_valid);
  always @(*) begin
    execute_ctrl2_down_MUL_SRC1_lane0 = _zz_execute_ctrl2_down_MUL_SRC1_lane0;
    if(execute_ctrl2_down_FpuMulPlugin_SEL_lane0) begin
      execute_ctrl2_down_MUL_SRC1_lane0 = {1'd0, FpuMulPlugin_logic_mulCmd_m1};
    end
  end

  always @(*) begin
    execute_ctrl2_down_MUL_SRC2_lane0 = _zz_execute_ctrl2_down_MUL_SRC2_lane0;
    if(execute_ctrl2_down_FpuMulPlugin_SEL_lane0) begin
      execute_ctrl2_down_MUL_SRC2_lane0 = {1'd0, FpuMulPlugin_logic_mulCmd_m2};
    end
  end

  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[33 : 17] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[33 : 17]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[50 : 34] * execute_ctrl2_down_MUL_SRC2_lane0[50 : 34]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[33 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[50 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[50 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6[60 : 51] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0[9 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[43 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0[36 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1[43 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[53 : 10];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2[43 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[53 : 10];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3[43 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0[36 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[6 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0[33 : 27];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[40 : 7] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4[43 : 41] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0[2 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5[23 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0[33 : 10];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5[43 : 24] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0[19 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6 = 44'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6[23 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0[33 : 10];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6[43 : 24] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0[19 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0[39 : 37];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_1[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0[56 : 54];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_2[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0[56 : 54];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_3[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0[39 : 37];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_4[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0[5 : 3];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_5[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0[22 : 20];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_6[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0[22 : 20];
  end

  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_14);
  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_14);
  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_7 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0_14);
  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = 111'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 0] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[63 : 0];
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[110 : 105] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0[5 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1 = 111'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1[107 : 61] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[46 : 0];
  end

  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = (_zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 + _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1);
  assign early0_MulPlugin_logic_formatBus_valid = execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  assign early0_MulPlugin_logic_formatBus_payload = (execute_ctrl4_down_MulPlugin_HIGH_lane0 ? execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 32] : execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[31 : 0]);
  assign io_cmd_fire = (early0_DivPlugin_logic_processing_div_io_cmd_valid && early0_DivPlugin_logic_processing_div_io_cmd_ready);
  always @(*) begin
    early0_DivPlugin_logic_processing_request = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_DivPlugin_SEL_lane0);
    if(when_FpuDivPlugin_l68) begin
      early0_DivPlugin_logic_processing_request = 1'b1;
    end
  end

  always @(*) begin
    early0_DivPlugin_logic_processing_a = {32'd0, execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0};
    if(when_FpuDivPlugin_l68) begin
      early0_DivPlugin_logic_processing_a = {11'd0, _zz_early0_DivPlugin_logic_processing_a};
    end
  end

  always @(*) begin
    early0_DivPlugin_logic_processing_b = {32'd0, execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0};
    if(when_FpuDivPlugin_l68) begin
      early0_DivPlugin_logic_processing_b = {11'd0, _zz_early0_DivPlugin_logic_processing_b};
    end
  end

  assign early0_DivPlugin_logic_processing_div_io_cmd_valid = (early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_cmdSent));
  always @(*) begin
    early0_DivPlugin_logic_processing_div_io_cmd_payload_normalized = 1'b0;
    if(when_FpuDivPlugin_l68) begin
      early0_DivPlugin_logic_processing_div_io_cmd_payload_normalized = 1'b1;
    end
  end

  always @(*) begin
    early0_DivPlugin_logic_processing_div_io_cmd_payload_iterations = 5'bxxxxx;
    if(when_FpuDivPlugin_l68) begin
      early0_DivPlugin_logic_processing_div_io_cmd_payload_iterations = 5'h1c;
    end
  end

  assign early0_DivPlugin_logic_processing_freeze = ((early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_div_io_rsp_valid)) && (! early0_DivPlugin_logic_processing_unscheduleRequest));
  assign early0_DivPlugin_logic_processing_selected = (execute_ctrl2_down_DivPlugin_REM_lane0 ? _zz_early0_DivPlugin_logic_processing_selected : _zz_early0_DivPlugin_logic_processing_selected_1);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = early0_DivPlugin_logic_processing_selected;
  assign execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  assign early0_DivPlugin_logic_formatBus_valid = execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  assign early0_DivPlugin_logic_formatBus_payload = execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  assign early0_EnvPlugin_logic_exe_privilege = PrivilegedPlugin_logic_harts_0_privilege;
  assign early0_EnvPlugin_logic_exe_xretPriv = execute_ctrl2_down_Decode_UOP_lane0[29 : 28];
  always @(*) begin
    early0_EnvPlugin_logic_exe_commit = 1'b0;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_exe_commit = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_retKo = 1'b0;
  assign early0_EnvPlugin_logic_exe_vmaKo = 1'b0;
  assign when_EnvPlugin_l86 = ((early0_EnvPlugin_logic_exe_xretPriv <= PrivilegedPlugin_logic_harts_0_privilege) && (! early0_EnvPlugin_logic_exe_retKo));
  assign when_EnvPlugin_l95 = ((early0_EnvPlugin_logic_exe_privilege == 2'b11) || ((! PrivilegedPlugin_logic_harts_0_m_status_tw) && (1'b1 || (early0_EnvPlugin_logic_exe_privilege == 2'b01))));
  assign when_EnvPlugin_l119 = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_EnvPlugin_SEL_lane0);
  assign when_EnvPlugin_l123 = (! early0_EnvPlugin_logic_exe_commit);
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_PC_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early0_BranchPlugin_pcCalc_target_b = {{11{_zz_early0_BranchPlugin_pcCalc_target_b[20]}}, _zz_early0_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_b = {{20{_zz_early0_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early0_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_b = {{19{_zz_early0_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early0_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early0_BranchPlugin_pcCalc_slices = ({1'b0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} + {1'b0,1'b1});
  always @(*) begin
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0] = 1'b0;
  end

  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0);
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early1_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1;
      end
      default : begin
        early1_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_PC_lane1;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early1_BranchPlugin_pcCalc_target_b = {{11{_zz_early1_BranchPlugin_pcCalc_target_b[20]}}, _zz_early1_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early1_BranchPlugin_pcCalc_target_b = {{20{_zz_early1_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early1_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early1_BranchPlugin_pcCalc_target_b = {{19{_zz_early1_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early1_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early1_BranchPlugin_pcCalc_slices = ({1'b0,execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1} + {1'b0,1'b1});
  always @(*) begin
    execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
    execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0] = 1'b0;
  end

  assign execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = (execute_ctrl2_down_PC_lane1 + _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = (execute_ctrl2_down_PC_lane1 + _zz_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1);
  assign AlignerPlugin_logic_maskGen_frontMasks_0 = 4'b1111;
  assign AlignerPlugin_logic_maskGen_frontMasks_1 = 4'b1110;
  assign AlignerPlugin_logic_maskGen_frontMasks_2 = 4'b1100;
  assign AlignerPlugin_logic_maskGen_frontMasks_3 = 4'b1000;
  assign AlignerPlugin_logic_maskGen_backMasks_0 = 4'b0001;
  assign AlignerPlugin_logic_maskGen_backMasks_1 = 4'b0011;
  assign AlignerPlugin_logic_maskGen_backMasks_2 = 4'b0111;
  assign AlignerPlugin_logic_maskGen_backMasks_3 = 4'b1111;
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = (_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & ((! fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? 4'b1111 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2));
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = ((fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST : 4'b0000);
  assign AlignerPlugin_logic_slicesInstructions_0 = {AlignerPlugin_logic_slices_data_1,AlignerPlugin_logic_slices_data_0};
  assign AlignerPlugin_logic_slicesInstructions_1 = {AlignerPlugin_logic_slices_data_2,AlignerPlugin_logic_slices_data_1};
  assign AlignerPlugin_logic_slicesInstructions_2 = {AlignerPlugin_logic_slices_data_3,AlignerPlugin_logic_slices_data_2};
  assign AlignerPlugin_logic_slicesInstructions_3 = {AlignerPlugin_logic_slices_data_4,AlignerPlugin_logic_slices_data_3};
  assign AlignerPlugin_logic_slicesInstructions_4 = {AlignerPlugin_logic_slices_data_5,AlignerPlugin_logic_slices_data_4};
  assign AlignerPlugin_logic_slicesInstructions_5 = {AlignerPlugin_logic_slices_data_6,AlignerPlugin_logic_slices_data_5};
  assign AlignerPlugin_logic_slicesInstructions_6 = {AlignerPlugin_logic_slices_data_7,AlignerPlugin_logic_slices_data_6};
  assign AlignerPlugin_logic_slicesInstructions_7 = {16'd0, AlignerPlugin_logic_slices_data_7};
  always @(*) begin
    AlignerPlugin_logic_scanners_0_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_0_usageMask[0] = AlignerPlugin_logic_scanners_0_checker_0_required;
    AlignerPlugin_logic_scanners_0_usageMask[1] = AlignerPlugin_logic_scanners_0_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_0_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_0_checker_0_last = (AlignerPlugin_logic_slices_data_0[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_0_redo = ((AlignerPlugin_logic_scanners_0_checker_0_required && AlignerPlugin_logic_slices_last[0]) && (! AlignerPlugin_logic_scanners_0_checker_0_last));
  assign AlignerPlugin_logic_scanners_0_checker_0_present = AlignerPlugin_logic_slices_mask[0];
  assign AlignerPlugin_logic_scanners_0_checker_0_valid = AlignerPlugin_logic_scanners_0_checker_0_present;
  assign AlignerPlugin_logic_scanners_0_checker_1_required = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_last = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_redo = ((AlignerPlugin_logic_scanners_0_checker_1_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_0_checker_1_last));
  assign AlignerPlugin_logic_scanners_0_checker_1_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_0_checker_1_valid = (AlignerPlugin_logic_scanners_0_checker_1_present || (! AlignerPlugin_logic_scanners_0_checker_1_required));
  assign AlignerPlugin_logic_scanners_0_redo = (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo});
  assign AlignerPlugin_logic_scanners_0_valid = (AlignerPlugin_logic_scanners_0_checker_0_valid && ((&AlignerPlugin_logic_scanners_0_checker_1_valid) || (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_1_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_1_usageMask[1] = AlignerPlugin_logic_scanners_1_checker_0_required;
    AlignerPlugin_logic_scanners_1_usageMask[2] = AlignerPlugin_logic_scanners_1_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_1_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_1_checker_0_last = (AlignerPlugin_logic_slices_data_1[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_0_redo = ((AlignerPlugin_logic_scanners_1_checker_0_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_1_checker_0_last));
  assign AlignerPlugin_logic_scanners_1_checker_0_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_1_checker_0_valid = AlignerPlugin_logic_scanners_1_checker_0_present;
  assign AlignerPlugin_logic_scanners_1_checker_1_required = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_last = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_redo = ((AlignerPlugin_logic_scanners_1_checker_1_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_1_checker_1_last));
  assign AlignerPlugin_logic_scanners_1_checker_1_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_1_checker_1_valid = (AlignerPlugin_logic_scanners_1_checker_1_present || (! AlignerPlugin_logic_scanners_1_checker_1_required));
  assign AlignerPlugin_logic_scanners_1_redo = (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo});
  assign AlignerPlugin_logic_scanners_1_valid = (AlignerPlugin_logic_scanners_1_checker_0_valid && ((&AlignerPlugin_logic_scanners_1_checker_1_valid) || (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_2_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_2_usageMask[2] = AlignerPlugin_logic_scanners_2_checker_0_required;
    AlignerPlugin_logic_scanners_2_usageMask[3] = AlignerPlugin_logic_scanners_2_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_2_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_2_checker_0_last = (AlignerPlugin_logic_slices_data_2[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_0_redo = ((AlignerPlugin_logic_scanners_2_checker_0_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_2_checker_0_last));
  assign AlignerPlugin_logic_scanners_2_checker_0_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_2_checker_0_valid = AlignerPlugin_logic_scanners_2_checker_0_present;
  assign AlignerPlugin_logic_scanners_2_checker_1_required = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_last = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_redo = ((AlignerPlugin_logic_scanners_2_checker_1_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_2_checker_1_last));
  assign AlignerPlugin_logic_scanners_2_checker_1_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_2_checker_1_valid = (AlignerPlugin_logic_scanners_2_checker_1_present || (! AlignerPlugin_logic_scanners_2_checker_1_required));
  assign AlignerPlugin_logic_scanners_2_redo = (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo});
  assign AlignerPlugin_logic_scanners_2_valid = (AlignerPlugin_logic_scanners_2_checker_0_valid && ((&AlignerPlugin_logic_scanners_2_checker_1_valid) || (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_3_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_3_usageMask[3] = AlignerPlugin_logic_scanners_3_checker_0_required;
    AlignerPlugin_logic_scanners_3_usageMask[4] = AlignerPlugin_logic_scanners_3_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_3_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_3_checker_0_last = (AlignerPlugin_logic_slices_data_3[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_0_redo = ((AlignerPlugin_logic_scanners_3_checker_0_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_3_checker_0_last));
  assign AlignerPlugin_logic_scanners_3_checker_0_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_3_checker_0_valid = AlignerPlugin_logic_scanners_3_checker_0_present;
  assign AlignerPlugin_logic_scanners_3_checker_1_required = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_last = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_redo = ((AlignerPlugin_logic_scanners_3_checker_1_required && AlignerPlugin_logic_slices_last[4]) && (! AlignerPlugin_logic_scanners_3_checker_1_last));
  assign AlignerPlugin_logic_scanners_3_checker_1_present = AlignerPlugin_logic_slices_mask[4];
  assign AlignerPlugin_logic_scanners_3_checker_1_valid = (AlignerPlugin_logic_scanners_3_checker_1_present || (! AlignerPlugin_logic_scanners_3_checker_1_required));
  assign AlignerPlugin_logic_scanners_3_redo = (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo});
  assign AlignerPlugin_logic_scanners_3_valid = (AlignerPlugin_logic_scanners_3_checker_0_valid && ((&AlignerPlugin_logic_scanners_3_checker_1_valid) || (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_4_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_4_usageMask[4] = AlignerPlugin_logic_scanners_4_checker_0_required;
    AlignerPlugin_logic_scanners_4_usageMask[5] = AlignerPlugin_logic_scanners_4_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_4_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_4_checker_0_last = (AlignerPlugin_logic_slices_data_4[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_0_redo = ((AlignerPlugin_logic_scanners_4_checker_0_required && AlignerPlugin_logic_slices_last[4]) && (! AlignerPlugin_logic_scanners_4_checker_0_last));
  assign AlignerPlugin_logic_scanners_4_checker_0_present = AlignerPlugin_logic_slices_mask[4];
  assign AlignerPlugin_logic_scanners_4_checker_0_valid = AlignerPlugin_logic_scanners_4_checker_0_present;
  assign AlignerPlugin_logic_scanners_4_checker_1_required = (AlignerPlugin_logic_slices_data_4[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_1_last = (AlignerPlugin_logic_slices_data_4[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_1_redo = ((AlignerPlugin_logic_scanners_4_checker_1_required && AlignerPlugin_logic_slices_last[5]) && (! AlignerPlugin_logic_scanners_4_checker_1_last));
  assign AlignerPlugin_logic_scanners_4_checker_1_present = AlignerPlugin_logic_slices_mask[5];
  assign AlignerPlugin_logic_scanners_4_checker_1_valid = (AlignerPlugin_logic_scanners_4_checker_1_present || (! AlignerPlugin_logic_scanners_4_checker_1_required));
  assign AlignerPlugin_logic_scanners_4_redo = (|{AlignerPlugin_logic_scanners_4_checker_1_redo,AlignerPlugin_logic_scanners_4_checker_0_redo});
  assign AlignerPlugin_logic_scanners_4_valid = (AlignerPlugin_logic_scanners_4_checker_0_valid && ((&AlignerPlugin_logic_scanners_4_checker_1_valid) || (|{AlignerPlugin_logic_scanners_4_checker_1_redo,AlignerPlugin_logic_scanners_4_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_5_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_5_usageMask[5] = AlignerPlugin_logic_scanners_5_checker_0_required;
    AlignerPlugin_logic_scanners_5_usageMask[6] = AlignerPlugin_logic_scanners_5_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_5_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_5_checker_0_last = (AlignerPlugin_logic_slices_data_5[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_0_redo = ((AlignerPlugin_logic_scanners_5_checker_0_required && AlignerPlugin_logic_slices_last[5]) && (! AlignerPlugin_logic_scanners_5_checker_0_last));
  assign AlignerPlugin_logic_scanners_5_checker_0_present = AlignerPlugin_logic_slices_mask[5];
  assign AlignerPlugin_logic_scanners_5_checker_0_valid = AlignerPlugin_logic_scanners_5_checker_0_present;
  assign AlignerPlugin_logic_scanners_5_checker_1_required = (AlignerPlugin_logic_slices_data_5[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_1_last = (AlignerPlugin_logic_slices_data_5[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_1_redo = ((AlignerPlugin_logic_scanners_5_checker_1_required && AlignerPlugin_logic_slices_last[6]) && (! AlignerPlugin_logic_scanners_5_checker_1_last));
  assign AlignerPlugin_logic_scanners_5_checker_1_present = AlignerPlugin_logic_slices_mask[6];
  assign AlignerPlugin_logic_scanners_5_checker_1_valid = (AlignerPlugin_logic_scanners_5_checker_1_present || (! AlignerPlugin_logic_scanners_5_checker_1_required));
  assign AlignerPlugin_logic_scanners_5_redo = (|{AlignerPlugin_logic_scanners_5_checker_1_redo,AlignerPlugin_logic_scanners_5_checker_0_redo});
  assign AlignerPlugin_logic_scanners_5_valid = (AlignerPlugin_logic_scanners_5_checker_0_valid && ((&AlignerPlugin_logic_scanners_5_checker_1_valid) || (|{AlignerPlugin_logic_scanners_5_checker_1_redo,AlignerPlugin_logic_scanners_5_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_6_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_6_usageMask[6] = AlignerPlugin_logic_scanners_6_checker_0_required;
    AlignerPlugin_logic_scanners_6_usageMask[7] = AlignerPlugin_logic_scanners_6_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_6_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_6_checker_0_last = (AlignerPlugin_logic_slices_data_6[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_0_redo = ((AlignerPlugin_logic_scanners_6_checker_0_required && AlignerPlugin_logic_slices_last[6]) && (! AlignerPlugin_logic_scanners_6_checker_0_last));
  assign AlignerPlugin_logic_scanners_6_checker_0_present = AlignerPlugin_logic_slices_mask[6];
  assign AlignerPlugin_logic_scanners_6_checker_0_valid = AlignerPlugin_logic_scanners_6_checker_0_present;
  assign AlignerPlugin_logic_scanners_6_checker_1_required = (AlignerPlugin_logic_slices_data_6[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_1_last = (AlignerPlugin_logic_slices_data_6[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_1_redo = ((AlignerPlugin_logic_scanners_6_checker_1_required && AlignerPlugin_logic_slices_last[7]) && (! AlignerPlugin_logic_scanners_6_checker_1_last));
  assign AlignerPlugin_logic_scanners_6_checker_1_present = AlignerPlugin_logic_slices_mask[7];
  assign AlignerPlugin_logic_scanners_6_checker_1_valid = (AlignerPlugin_logic_scanners_6_checker_1_present || (! AlignerPlugin_logic_scanners_6_checker_1_required));
  assign AlignerPlugin_logic_scanners_6_redo = (|{AlignerPlugin_logic_scanners_6_checker_1_redo,AlignerPlugin_logic_scanners_6_checker_0_redo});
  assign AlignerPlugin_logic_scanners_6_valid = (AlignerPlugin_logic_scanners_6_checker_0_valid && ((&AlignerPlugin_logic_scanners_6_checker_1_valid) || (|{AlignerPlugin_logic_scanners_6_checker_1_redo,AlignerPlugin_logic_scanners_6_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_7_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_7_usageMask[7] = AlignerPlugin_logic_scanners_7_checker_0_required;
  end

  assign AlignerPlugin_logic_scanners_7_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_7_checker_0_last = (AlignerPlugin_logic_slices_data_7[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_0_redo = ((AlignerPlugin_logic_scanners_7_checker_0_required && AlignerPlugin_logic_slices_last[7]) && (! AlignerPlugin_logic_scanners_7_checker_0_last));
  assign AlignerPlugin_logic_scanners_7_checker_0_present = AlignerPlugin_logic_slices_mask[7];
  assign AlignerPlugin_logic_scanners_7_checker_0_valid = AlignerPlugin_logic_scanners_7_checker_0_present;
  assign AlignerPlugin_logic_scanners_7_checker_1_required = (AlignerPlugin_logic_slices_data_7[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_1_last = (AlignerPlugin_logic_slices_data_7[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_1_redo = 1'b0;
  assign AlignerPlugin_logic_scanners_7_checker_1_present = 1'b0;
  assign AlignerPlugin_logic_scanners_7_checker_1_valid = (AlignerPlugin_logic_scanners_7_checker_1_present || (! AlignerPlugin_logic_scanners_7_checker_1_required));
  assign AlignerPlugin_logic_scanners_7_redo = (|{AlignerPlugin_logic_scanners_7_checker_1_redo,AlignerPlugin_logic_scanners_7_checker_0_redo});
  assign AlignerPlugin_logic_scanners_7_valid = (AlignerPlugin_logic_scanners_7_checker_0_valid && ((&AlignerPlugin_logic_scanners_7_checker_1_valid) || (|{AlignerPlugin_logic_scanners_7_checker_1_redo,AlignerPlugin_logic_scanners_7_checker_0_redo})));
  assign AlignerPlugin_logic_usedMask_0 = 8'h0;
  assign AlignerPlugin_logic_extractors_0_first = 1'b1;
  assign AlignerPlugin_logic_extractors_0_usableMask = {(AlignerPlugin_logic_scanners_7_valid && (! AlignerPlugin_logic_usedMask_0[7])),{(AlignerPlugin_logic_scanners_6_valid && (! AlignerPlugin_logic_usedMask_0[6])),{(AlignerPlugin_logic_scanners_5_valid && (! AlignerPlugin_logic_usedMask_0[5])),{(AlignerPlugin_logic_scanners_4_valid && (! _zz_AlignerPlugin_logic_extractors_0_usableMask)),{(AlignerPlugin_logic_scanners_3_valid && _zz_AlignerPlugin_logic_extractors_0_usableMask_1),{_zz_AlignerPlugin_logic_extractors_0_usableMask_2,{_zz_AlignerPlugin_logic_extractors_0_usableMask_3,_zz_AlignerPlugin_logic_extractors_0_usableMask_4}}}}}}};
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0 = AlignerPlugin_logic_extractors_0_usableMask;
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_0 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[0];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_1 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[1];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_2 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[2];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_3 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[3];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_4 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[4];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_5 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[5];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_6 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[6];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_7 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[7];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[0] = (AlignerPlugin_logic_extractors_0_usableMask_bools_0 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[1] = (AlignerPlugin_logic_extractors_0_usableMask_bools_1 && (! AlignerPlugin_logic_extractors_0_usableMask_bools_0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[2] = (AlignerPlugin_logic_extractors_0_usableMask_bools_2 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[3] = (AlignerPlugin_logic_extractors_0_usableMask_bools_3 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[4] = (AlignerPlugin_logic_extractors_0_usableMask_bools_4 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[5] = (AlignerPlugin_logic_extractors_0_usableMask_bools_5 && (! (AlignerPlugin_logic_extractors_0_usableMask_bools_4 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[6] = (AlignerPlugin_logic_extractors_0_usableMask_bools_6 && (! (AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[7] = (AlignerPlugin_logic_extractors_0_usableMask_bools_7 && (! (AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
  end

  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_2,{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0}});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_3,{AlignerPlugin_logic_extractors_0_usableMask_bools_2,{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0}}});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_5,AlignerPlugin_logic_extractors_0_usableMask_bools_4});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_6,{AlignerPlugin_logic_extractors_0_usableMask_bools_5,AlignerPlugin_logic_extractors_0_usableMask_bools_4}});
  assign AlignerPlugin_logic_extractors_0_slicesOh = _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  assign _zz_AlignerPlugin_logic_extractors_0_redo = AlignerPlugin_logic_extractors_0_slicesOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_1 = AlignerPlugin_logic_extractors_0_slicesOh[1];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_2 = AlignerPlugin_logic_extractors_0_slicesOh[2];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_3 = AlignerPlugin_logic_extractors_0_slicesOh[3];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_4 = AlignerPlugin_logic_extractors_0_slicesOh[4];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_5 = AlignerPlugin_logic_extractors_0_slicesOh[5];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_6 = AlignerPlugin_logic_extractors_0_slicesOh[6];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_7 = AlignerPlugin_logic_extractors_0_slicesOh[7];
  always @(*) begin
    AlignerPlugin_logic_extractors_0_redo = _zz_AlignerPlugin_logic_extractors_0_redo_8[0];
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_0_localMask = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? {_zz_AlignerPlugin_logic_extractors_0_localMask,_zz_AlignerPlugin_logic_extractors_0_localMask_1} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_2,_zz_AlignerPlugin_logic_extractors_0_localMask_3} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_4,_zz_AlignerPlugin_logic_extractors_0_localMask_5} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_6,_zz_AlignerPlugin_logic_extractors_0_localMask_7} : 2'b00))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_8,_zz_AlignerPlugin_logic_extractors_0_localMask_9} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_10,_zz_AlignerPlugin_logic_extractors_0_localMask_11} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_12,_zz_AlignerPlugin_logic_extractors_0_localMask_13} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_14,_zz_AlignerPlugin_logic_extractors_0_localMask_15} : 2'b00))));
  assign AlignerPlugin_logic_extractors_0_usageMask = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? AlignerPlugin_logic_scanners_0_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? AlignerPlugin_logic_scanners_1_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? AlignerPlugin_logic_scanners_2_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? AlignerPlugin_logic_scanners_3_usageMask : 8'h0))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? AlignerPlugin_logic_scanners_4_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? AlignerPlugin_logic_scanners_5_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? AlignerPlugin_logic_scanners_6_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? AlignerPlugin_logic_scanners_7_usageMask : 8'h0))));
  assign AlignerPlugin_logic_usedMask_1 = (AlignerPlugin_logic_usedMask_0 | AlignerPlugin_logic_extractors_0_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_0_valid = (|AlignerPlugin_logic_extractors_0_slicesOh);
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_valid = 1'b0;
    end
    if(when_AlignerPlugin_l240) begin
      if(when_AlignerPlugin_l241) begin
        AlignerPlugin_logic_extractors_0_valid = 1'b0;
      end
    end
  end

  assign when_AlignerPlugin_l160 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_0_first)));
  assign AlignerPlugin_logic_extractors_1_first = 1'b0;
  assign AlignerPlugin_logic_extractors_1_usableMask = {(AlignerPlugin_logic_scanners_7_valid && (! AlignerPlugin_logic_usedMask_1[7])),{(AlignerPlugin_logic_scanners_6_valid && (! AlignerPlugin_logic_usedMask_1[6])),{(AlignerPlugin_logic_scanners_5_valid && (! AlignerPlugin_logic_usedMask_1[5])),{(AlignerPlugin_logic_scanners_4_valid && (! _zz_AlignerPlugin_logic_extractors_1_usableMask)),{(AlignerPlugin_logic_scanners_3_valid && _zz_AlignerPlugin_logic_extractors_1_usableMask_1),{_zz_AlignerPlugin_logic_extractors_1_usableMask_2,_zz_AlignerPlugin_logic_extractors_1_usableMask_3}}}}}};
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0 = AlignerPlugin_logic_extractors_1_usableMask;
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_0 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[0];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_1 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[1];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_2 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[2];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_3 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[3];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_4 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[4];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_5 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[5];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_6 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[6];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[0] = (AlignerPlugin_logic_extractors_1_usableMask_bools_0 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[1] = (AlignerPlugin_logic_extractors_1_usableMask_bools_1 && (! AlignerPlugin_logic_extractors_1_usableMask_bools_0));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[2] = (AlignerPlugin_logic_extractors_1_usableMask_bools_2 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[3] = (AlignerPlugin_logic_extractors_1_usableMask_bools_3 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[4] = (AlignerPlugin_logic_extractors_1_usableMask_bools_4 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[5] = (AlignerPlugin_logic_extractors_1_usableMask_bools_5 && (! (AlignerPlugin_logic_extractors_1_usableMask_bools_4 || AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[6] = (AlignerPlugin_logic_extractors_1_usableMask_bools_6 && (! (AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5 || AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3)));
  end

  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_2,{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0}});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_3,{AlignerPlugin_logic_extractors_1_usableMask_bools_2,{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0}}});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_5,AlignerPlugin_logic_extractors_1_usableMask_bools_4});
  assign AlignerPlugin_logic_extractors_1_slicesOh = _zz_AlignerPlugin_logic_extractors_1_slicesOh;
  assign _zz_AlignerPlugin_logic_extractors_1_redo = AlignerPlugin_logic_extractors_1_slicesOh[0];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_1 = AlignerPlugin_logic_extractors_1_slicesOh[1];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_2 = AlignerPlugin_logic_extractors_1_slicesOh[2];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_3 = AlignerPlugin_logic_extractors_1_slicesOh[3];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_4 = AlignerPlugin_logic_extractors_1_slicesOh[4];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_5 = AlignerPlugin_logic_extractors_1_slicesOh[5];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_6 = AlignerPlugin_logic_extractors_1_slicesOh[6];
  always @(*) begin
    AlignerPlugin_logic_extractors_1_redo = _zz_AlignerPlugin_logic_extractors_1_redo_7[0];
    if(when_AlignerPlugin_l160_1) begin
      AlignerPlugin_logic_extractors_1_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_1_localMask = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? {_zz_AlignerPlugin_logic_extractors_1_localMask,_zz_AlignerPlugin_logic_extractors_1_localMask_1} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_2,_zz_AlignerPlugin_logic_extractors_1_localMask_3} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_4,_zz_AlignerPlugin_logic_extractors_1_localMask_5} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_6,_zz_AlignerPlugin_logic_extractors_1_localMask_7} : 2'b00))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_8,_zz_AlignerPlugin_logic_extractors_1_localMask_9} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_10,_zz_AlignerPlugin_logic_extractors_1_localMask_11} : 2'b00)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? {AlignerPlugin_logic_scanners_7_checker_1_required,AlignerPlugin_logic_scanners_7_checker_0_required} : 2'b00)));
  assign AlignerPlugin_logic_extractors_1_usageMask = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? AlignerPlugin_logic_scanners_1_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? AlignerPlugin_logic_scanners_2_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? AlignerPlugin_logic_scanners_3_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? AlignerPlugin_logic_scanners_4_usageMask : 8'h0))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? AlignerPlugin_logic_scanners_5_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? AlignerPlugin_logic_scanners_6_usageMask : 8'h0)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? AlignerPlugin_logic_scanners_7_usageMask : 8'h0)));
  assign AlignerPlugin_logic_usedMask_2 = (AlignerPlugin_logic_usedMask_1 | AlignerPlugin_logic_extractors_1_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_1_valid = (|AlignerPlugin_logic_extractors_1_slicesOh);
    if(when_AlignerPlugin_l160_1) begin
      AlignerPlugin_logic_extractors_1_valid = 1'b0;
    end
    if(when_AlignerPlugin_l240) begin
      if(when_AlignerPlugin_l241_1) begin
        AlignerPlugin_logic_extractors_1_valid = 1'b0;
      end
    end
  end

  assign when_AlignerPlugin_l160_1 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_1_first)));
  assign when_AlignerPlugin_l171 = (decode_ctrls_0_up_isFiring && 1'b1);
  assign AlignerPlugin_logic_feeder_lanes_0_valid = AlignerPlugin_logic_extractors_0_valid;
  assign decode_ctrls_0_up_LANE_SEL_0 = AlignerPlugin_logic_feeder_lanes_0_valid;
  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = 1'b0;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_0_isRvc = (AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0] != 2'b11);
  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(switch_Rvc_l55)
      5'h0 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{{2'b00,AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00},5'h02},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h13};
      end
      5'h01 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h07};
      end
      5'h02 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h03};
      end
      5'h03 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h07};
      end
      5'h05 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[4 : 0]},7'h27};
      end
      5'h06 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[4 : 0]},7'h23};
      end
      5'h07 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[4 : 0]},7'h27};
      end
      5'h08 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h09 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[20],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[11]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20},7'h6f};
      end
      5'h0a : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,5'h0},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h0b : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h02) ? {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},4'b0000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13} : {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26[31 : 12],AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h37});
      end
      5'h0c : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27;
      end
      5'h0d : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[20],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[11]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},7'h6f};
      end
      5'h0e : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h0f : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b001},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h10 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{6'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b001},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h11 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{3'b000,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b011},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h07};
      end
      5'h12 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h03};
      end
      5'h13 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h07};
      end
      5'h14 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 2] == 11'h400) ? 32'h00100073 : ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) ? {{{{12'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19)},7'h67} : {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32},(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33 ? _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19)},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h33}));
      end
      5'h15 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36[4 : 0]},7'h27};
      end
      5'h16 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_37[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_38[4 : 0]},7'h23};
      end
      5'h17 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_39[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_40[4 : 0]},7'h27};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b0;
    case(switch_Rvc_l55)
      5'h0 : begin
        if(when_Rvc_l59) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h01 : begin
      end
      5'h02 : begin
      end
      5'h03 : begin
      end
      5'h05 : begin
      end
      5'h06 : begin
      end
      5'h07 : begin
      end
      5'h08 : begin
      end
      5'h09 : begin
      end
      5'h0a : begin
      end
      5'h0b : begin
        if(when_Rvc_l80) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0c : begin
      end
      5'h0d : begin
      end
      5'h0e : begin
      end
      5'h0f : begin
      end
      5'h10 : begin
      end
      5'h11 : begin
      end
      5'h12 : begin
        if(when_Rvc_l101) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h13 : begin
      end
      5'h14 : begin
        if(when_Rvc_l114) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h15 : begin
      end
      5'h16 : begin
      end
      5'h17 : begin
      end
      default : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
      end
    endcase
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1 = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 2]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2 = {{{{5'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[4 : 0] = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7,AlignerPlugin_logic_extractors_0_ctx_instruction[8]},AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},AlignerPlugin_logic_extractors_0_ctx_instruction[7]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[14] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[13] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[12] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14,AlignerPlugin_logic_extractors_0_ctx_instruction[8]},AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},AlignerPlugin_logic_extractors_0_ctx_instruction[7]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18 = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19 = 5'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20 = 5'h01;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21 = 5'h02;
  assign switch_Rvc_l55 = {AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0],AlignerPlugin_logic_extractors_0_ctx_instruction[15 : 13]};
  assign when_Rvc_l59 = (AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 5] == 8'h0);
  assign when_Rvc_l80 = ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 = {{{{_zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b101},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
  assign when_Rvc_l101 = (AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l114 = (((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0)) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = AlignerPlugin_logic_extractors_0_localMask;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[1]};
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[0];
  always @(*) begin
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[0] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 && (! 1'b0));
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[1] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[1] && (! _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2));
  end

  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5[1];
  assign decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  assign decode_ctrls_0_up_PC_0 = AlignerPlugin_logic_extractors_0_ctx_pc;
  assign decode_ctrls_0_up_Decode_DOP_ID_0 = AlignerPlugin_logic_feeder_harts_0_dopId;
  assign decode_ctrls_0_up_Fetch_ID_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  assign decode_ctrls_0_up_Prediction_WORD_JUMPED_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  assign decode_ctrls_0_up_TRAP_0 = AlignerPlugin_logic_extractors_0_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice = (decode_ctrls_0_up_PC_0[2 : 1] + _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice);
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction = (decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 <= AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0 = (decode_ctrls_0_up_Prediction_WORD_JUMPED_0 && AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  assign decode_ctrls_0_up_Prediction_ALIGN_REDO_0 = AlignerPlugin_logic_extractors_0_redo;
  assign AlignerPlugin_logic_feeder_lanes_1_valid = AlignerPlugin_logic_extractors_1_valid;
  assign decode_ctrls_0_up_LANE_SEL_1 = AlignerPlugin_logic_feeder_lanes_1_valid;
  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_1 = AlignerPlugin_logic_extractors_1_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_1 = AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1 = 1'b0;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1 = AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal;
    end
  end

  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1 = AlignerPlugin_logic_extractors_1_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_1_isRvc = (AlignerPlugin_logic_extractors_1_ctx_instruction[1 : 0] != 2'b11);
  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(switch_Rvc_l55_1)
      5'h0 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{{2'b00,AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},2'b00},5'h02},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h13};
      end
      5'h01 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h07};
      end
      5'h02 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h03};
      end
      5'h03 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h07};
      end
      5'h05 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3[4 : 0]},7'h27};
      end
      5'h06 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[4 : 0]},7'h23};
      end
      5'h07 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[4 : 0]},7'h27};
      end
      5'h08 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h09 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[20],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[11]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20},7'h6f};
      end
      5'h0a : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,5'h0},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h0b : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h02) ? {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},4'b0000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13} : {{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26[31 : 12],AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h37});
      end
      5'h0c : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27;
      end
      5'h0d : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[20],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[11]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},7'h6f};
      end
      5'h0e : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h0f : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b001},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h10 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{6'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b001},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h11 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{3'b000,AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b011},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h07};
      end
      5'h12 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h03};
      end
      5'h13 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h07};
      end
      5'h14 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 2] == 11'h400) ? 32'h00100073 : ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0) ? {{{{12'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},(AlignerPlugin_logic_extractors_1_ctx_instruction[12] ? _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19)},7'h67} : {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32},(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33 ? _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19)},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h33}));
      end
      5'h15 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35[11 : 5],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36[4 : 0]},7'h27};
      end
      5'h16 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_37[11 : 5],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_38[4 : 0]},7'h23};
      end
      5'h17 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_39[11 : 5],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_40[4 : 0]},7'h27};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b0;
    case(switch_Rvc_l55_1)
      5'h0 : begin
        if(when_Rvc_l59_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h01 : begin
      end
      5'h02 : begin
      end
      5'h03 : begin
      end
      5'h05 : begin
      end
      5'h06 : begin
      end
      5'h07 : begin
      end
      5'h08 : begin
      end
      5'h09 : begin
      end
      5'h0a : begin
      end
      5'h0b : begin
        if(when_Rvc_l80_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0c : begin
      end
      5'h0d : begin
      end
      5'h0e : begin
      end
      5'h0f : begin
      end
      5'h10 : begin
      end
      5'h11 : begin
      end
      5'h12 : begin
        if(when_Rvc_l101_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h13 : begin
      end
      5'h14 : begin
        if(when_Rvc_l114_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h15 : begin
      end
      5'h16 : begin
      end
      5'h17 : begin
      end
      default : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
      end
    endcase
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {2'b01,AlignerPlugin_logic_extractors_1_ctx_instruction[9 : 7]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1 = {2'b01,AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 2]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2 = {{{{5'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[5]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[11] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[10] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[4 : 0] = AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2];
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7,AlignerPlugin_logic_extractors_1_ctx_instruction[8]},AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},AlignerPlugin_logic_extractors_1_ctx_instruction[7]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[14] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[13] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[12] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[11] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[10] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14,AlignerPlugin_logic_extractors_1_ctx_instruction[8]},AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},AlignerPlugin_logic_extractors_1_ctx_instruction[7]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18 = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 10]},AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19 = 5'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20 = 5'h01;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21 = 5'h02;
  assign switch_Rvc_l55_1 = {AlignerPlugin_logic_extractors_1_ctx_instruction[1 : 0],AlignerPlugin_logic_extractors_1_ctx_instruction[15 : 13]};
  assign when_Rvc_l59_1 = (AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 5] == 8'h0);
  assign when_Rvc_l80_1 = ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0) && (AlignerPlugin_logic_extractors_1_ctx_instruction[12] == 1'b0));
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 = {{{{_zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b101},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},7'h13};
  assign when_Rvc_l101_1 = (AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l114_1 = (((AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h0) && (AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0)) && (AlignerPlugin_logic_extractors_1_ctx_instruction[12] == 1'b0));
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1 = AlignerPlugin_logic_extractors_1_localMask;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1 = {_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1[0],_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1[1]};
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1[0];
  always @(*) begin
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3[0] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2 && (! 1'b0));
    _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3[1] = (_zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1[1] && (! _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2));
  end

  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3;
  assign _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5 = _zz__zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5[1];
  assign decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1 = _zz_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  assign decode_ctrls_0_up_PC_1 = AlignerPlugin_logic_extractors_1_ctx_pc;
  assign decode_ctrls_0_up_Decode_DOP_ID_1 = (decode_ctrls_0_down_Decode_DOP_ID_0 + _zz_decode_ctrls_0_up_Decode_DOP_ID_1);
  assign decode_ctrls_0_up_Fetch_ID_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC;
  assign decode_ctrls_0_up_Prediction_WORD_JUMPED_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE;
  assign decode_ctrls_0_up_TRAP_1 = AlignerPlugin_logic_extractors_1_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice = (decode_ctrls_0_up_PC_1[2 : 1] + _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice);
  assign AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction = (decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1 <= AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1 = (decode_ctrls_0_up_Prediction_WORD_JUMPED_1 && AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1 = decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1 = decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1 = decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1;
  assign decode_ctrls_0_up_Prediction_ALIGN_REDO_1 = AlignerPlugin_logic_extractors_1_redo;
  assign decode_ctrls_0_up_valid = (|{AlignerPlugin_logic_feeder_lanes_1_valid,AlignerPlugin_logic_feeder_lanes_0_valid});
  assign _zz_AlignerPlugin_logic_slices_data_0 = {fetch_logic_ctrls_2_down_Fetch_WORD,AlignerPlugin_logic_buffer_data};
  assign AlignerPlugin_logic_slices_data_0 = _zz_AlignerPlugin_logic_slices_data_0[15 : 0];
  assign AlignerPlugin_logic_slices_data_1 = _zz_AlignerPlugin_logic_slices_data_0[31 : 16];
  assign AlignerPlugin_logic_slices_data_2 = _zz_AlignerPlugin_logic_slices_data_0[47 : 32];
  assign AlignerPlugin_logic_slices_data_3 = _zz_AlignerPlugin_logic_slices_data_0[63 : 48];
  assign AlignerPlugin_logic_slices_data_4 = _zz_AlignerPlugin_logic_slices_data_0[79 : 64];
  assign AlignerPlugin_logic_slices_data_5 = _zz_AlignerPlugin_logic_slices_data_0[95 : 80];
  assign AlignerPlugin_logic_slices_data_6 = _zz_AlignerPlugin_logic_slices_data_0[111 : 96];
  assign AlignerPlugin_logic_slices_data_7 = _zz_AlignerPlugin_logic_slices_data_0[127 : 112];
  assign AlignerPlugin_logic_slices_mask = {(fetch_logic_ctrls_2_down_isValid ? fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK : 4'b0000),AlignerPlugin_logic_buffer_mask};
  assign AlignerPlugin_logic_slices_last = {fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST,AlignerPlugin_logic_buffer_last};
  assign when_AlignerPlugin_l240 = (! fetch_logic_ctrls_2_down_valid);
  assign when_AlignerPlugin_l241 = (AlignerPlugin_logic_extractors_0_usageMask[7 : 4] != 4'b0000);
  assign when_AlignerPlugin_l241_1 = (AlignerPlugin_logic_extractors_1_usageMask[7 : 4] != 4'b0000);
  assign AlignerPlugin_logic_buffer_downFire = (decode_ctrls_0_up_isReady || decode_ctrls_0_up_isCancel);
  assign AlignerPlugin_logic_buffer_usedMask = ((AlignerPlugin_logic_extractors_0_valid ? AlignerPlugin_logic_extractors_0_usageMask : 8'h0) | (AlignerPlugin_logic_extractors_1_valid ? AlignerPlugin_logic_extractors_1_usageMask : 8'h0));
  assign AlignerPlugin_logic_buffer_haltUp = ((|(AlignerPlugin_logic_buffer_mask & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[3 : 0] : 4'b0000)))) || AlignerPlugin_api_haltIt);
  assign fetch_logic_ctrls_2_down_ready = ((! fetch_logic_ctrls_2_down_valid) || (! AlignerPlugin_logic_buffer_haltUp));
  assign when_AlignerPlugin_l256 = ((fetch_logic_ctrls_2_down_isValid && fetch_logic_ctrls_2_down_isReady) && (! fetch_logic_ctrls_2_down_isCancel));
  assign _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0 = execute_ctrl2_down_Decode_UOP_lane0[14 : 12];
  assign _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1 = ((_zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0 == 3'b111) ? FpuCsrPlugin_api_rm : _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0);
  assign execute_ctrl2_down_FpuUtils_ROUNDING_lane0 = _zz_execute_ctrl2_down_FpuUtils_ROUNDING_lane0_1;
  assign when_FpuCsrPlugin_l61 = ((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_COMMIT_lane0) && execute_ctrl4_down_FpuCsrPlugin_DIRTY_lane0);
  assign execute_ctrl0_down_AguPlugin_SIZE_lane0 = execute_ctrl0_down_Decode_UOP_lane0[13 : 12];
  assign LsuPlugin_logic_storeBuffer_ops_full = (((LsuPlugin_logic_storeBuffer_ops_pushPtr ^ LsuPlugin_logic_storeBuffer_ops_freePtr) ^ 6'h20) == 6'h0);
  assign LsuPlugin_logic_storeBuffer_ops_occupancy = (LsuPlugin_logic_storeBuffer_ops_pushPtr - LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_0_valid = (LsuPlugin_logic_storeBuffer_ops_popPtr != LsuPlugin_logic_storeBuffer_ops_pushPtr);
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_0_SB_PTR = LsuPlugin_logic_storeBuffer_ops_popPtr;
  assign _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address = LsuPlugin_logic_storeBuffer_ops_popPtr;
  assign _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1 = LsuPlugin_logic_storeBuffer_ops_mem_spinal_port0;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address = _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1[31 : 0];
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_data = _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1[95 : 32];
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_size = _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1[97 : 96];
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_storeId = _zz_LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address_1[109 : 98];
  assign LsuPlugin_logic_storeBuffer_pop_valid = LsuPlugin_logic_storeBuffer_ops_pip_node_2_isValid;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_2_ready = LsuPlugin_logic_storeBuffer_pop_ready;
  assign LsuPlugin_logic_storeBuffer_pop_payload_op_address = LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_address;
  assign LsuPlugin_logic_storeBuffer_pop_payload_op_data = LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_data;
  assign LsuPlugin_logic_storeBuffer_pop_payload_op_size = LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_size;
  assign LsuPlugin_logic_storeBuffer_pop_payload_op_storeId = LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_storeId;
  assign LsuPlugin_logic_storeBuffer_pop_payload_ptr = LsuPlugin_logic_storeBuffer_ops_pip_node_2_SB_PTR;
  assign LsuPlugin_logic_storeBuffer_slotsFree = (|{(! LsuPlugin_logic_storeBuffer_slots_7_valid),{(! LsuPlugin_logic_storeBuffer_slots_6_valid),{(! LsuPlugin_logic_storeBuffer_slots_5_valid),{(! LsuPlugin_logic_storeBuffer_slots_4_valid),{(! LsuPlugin_logic_storeBuffer_slots_3_valid),{(! LsuPlugin_logic_storeBuffer_slots_2_valid),{(! LsuPlugin_logic_storeBuffer_slots_1_valid),(! LsuPlugin_logic_storeBuffer_slots_0_valid)}}}}}}});
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst = {(! LsuPlugin_logic_storeBuffer_slots_7_valid),{(! LsuPlugin_logic_storeBuffer_slots_6_valid),{(! LsuPlugin_logic_storeBuffer_slots_5_valid),{(! LsuPlugin_logic_storeBuffer_slots_4_valid),{(! LsuPlugin_logic_storeBuffer_slots_3_valid),{(! LsuPlugin_logic_storeBuffer_slots_2_valid),{(! LsuPlugin_logic_storeBuffer_slots_1_valid),(! LsuPlugin_logic_storeBuffer_slots_0_valid)}}}}}}};
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[0];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[1];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_3 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[2];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_4 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[3];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[4];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_6 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[5];
  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_7 = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[6];
  always @(*) begin
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[0] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1 && (! 1'b0));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[1] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2 && (! _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[2] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_3 && (! (|{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2,_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1})));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[3] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_4 && (! (|{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_3,{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2,_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1}})));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[4] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5 && (! _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[5] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_6 && (! (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5 || _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9)));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[6] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_7 && (! ((|{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_6,_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5}) || _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9)));
    _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8[7] = (_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst[7] && (! ((|{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_7,{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_6,_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_5}}) || _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9)));
  end

  assign _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_9 = (|{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_4,{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_3,{_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_2,_zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_1}}});
  assign LsuPlugin_logic_storeBuffer_slotsFreeFirst = _zz_LsuPlugin_logic_storeBuffer_slotsFreeFirst_8;
  assign when_LsuPlugin_l331 = (LsuPlugin_logic_storeBuffer_slotsFree && (LsuPlugin_logic_storeBuffer_ops_occupancy <= 6'h10));
  assign when_LsuPlugin_l259 = (|(LsuPlugin_logic_storeBuffer_waitL1_refill & (~ LsuL1_REFILL_BUSY)));
  assign LsuPlugin_logic_storeBuffer_empty = (&{(! LsuPlugin_logic_storeBuffer_slots_7_valid),{(! LsuPlugin_logic_storeBuffer_slots_6_valid),{(! LsuPlugin_logic_storeBuffer_slots_5_valid),{(! LsuPlugin_logic_storeBuffer_slots_4_valid),{(! LsuPlugin_logic_storeBuffer_slots_3_valid),{(! LsuPlugin_logic_storeBuffer_slots_2_valid),{(! LsuPlugin_logic_storeBuffer_slots_1_valid),(! LsuPlugin_logic_storeBuffer_slots_0_valid)}}}}}}});
  assign LsuPlugin_logic_flusher_wantExit = 1'b0;
  always @(*) begin
    LsuPlugin_logic_flusher_wantStart = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_SB_DRAIN : begin
      end
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
      end
      default : begin
        LsuPlugin_logic_flusher_wantStart = 1'b1;
      end
    endcase
  end

  assign LsuPlugin_logic_flusher_wantKill = 1'b0;
  assign TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready = LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_flusher_inflight = (|{(execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0),(execute_ctrl3_down_LsuL1_SEL_lane0 && execute_ctrl3_down_LsuL1_FLUSH_lane0)});
  always @(*) begin
    LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_SB_DRAIN : begin
      end
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l371) begin
          LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_api_lsuTriggerBus_load = execute_ctrl3_down_LsuL1_LOAD_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_store = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_virtual = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0 = 1'b0;
  assign execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = (execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 || execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0);
  assign LsuPlugin_logic_onAddress0_ls_prefetchOp = execute_ctrl2_down_Decode_UOP_lane0[24 : 20];
  assign LsuPlugin_logic_onAddress0_ls_port_valid = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_address = execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_size = execute_ctrl2_down_AguPlugin_SIZE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_load = execute_ctrl2_down_AguPlugin_LOAD_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_store = execute_ctrl2_down_AguPlugin_STORE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_atomic = execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_invalidate = 1'b0;
  always @(*) begin
    LsuPlugin_logic_onAddress0_ls_port_payload_op = LsuL1CmdOpcode_LSU;
    if(execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0) begin
      LsuPlugin_logic_onAddress0_ls_port_payload_op = LsuL1CmdOpcode_PREFETCH;
    end
  end

  assign LsuPlugin_logic_onAddress0_ls_port_fire = (LsuPlugin_logic_onAddress0_ls_port_valid && LsuPlugin_logic_onAddress0_ls_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_storeId = LsuPlugin_logic_onAddress0_ls_storeId;
  assign LsuPlugin_logic_onAddress0_flush_port_valid = ((LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD) && (! LsuPlugin_logic_flusher_cmdCounter[6]));
  assign LsuPlugin_logic_onAddress0_flush_port_payload_address = {19'd0, _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address};
  assign LsuPlugin_logic_onAddress0_flush_port_payload_size = 2'b00;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_op = LsuL1CmdOpcode_FLUSH;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_fire = (LsuPlugin_logic_onAddress0_flush_port_valid && LsuPlugin_logic_onAddress0_flush_port_ready);
  assign LsuPlugin_logic_onAddress0_sb_isHead = (LsuPlugin_logic_storeBuffer_pop_payload_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign LsuPlugin_logic_onAddress0_sb_flush = (LsuPlugin_logic_storeBuffer_waitL1_valid && (! LsuPlugin_logic_onAddress0_sb_isHead));
  assign LsuPlugin_logic_onAddress0_sb_port_valid = ((LsuPlugin_logic_storeBuffer_pop_valid && (! LsuPlugin_logic_storeBuffer_waitL1_valid)) && (! LsuPlugin_logic_onAddress0_sb_flush));
  assign LsuPlugin_logic_onAddress0_sb_port_payload_address = LsuPlugin_logic_storeBuffer_pop_payload_op_address;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_size = LsuPlugin_logic_storeBuffer_pop_payload_op_size;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_store = 1'b1;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_sb_port_payload_op = LsuL1CmdOpcode_STORE_BUFFER;
  assign LsuPlugin_logic_storeBuffer_pop_ready = (LsuPlugin_logic_onAddress0_sb_port_ready || LsuPlugin_logic_onAddress0_sb_flush);
  assign LsuPlugin_logic_onAddress0_sb_port_payload_storeId = LsuPlugin_logic_storeBuffer_pop_payload_op_storeId;
  assign LsuPlugin_logic_onAddress0_fromHp_port_valid = PrefetcherRptPlugin_io_valid;
  assign PrefetcherRptPlugin_io_ready = LsuPlugin_logic_onAddress0_fromHp_port_ready;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_op = LsuL1CmdOpcode_PREFETCH;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_address = PrefetcherRptPlugin_io_payload_address;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_store = PrefetcherRptPlugin_io_payload_unique;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_size = 2'b00;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_fromHp_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_ls_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_onAddress0_flush_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  assign LsuPlugin_logic_onAddress0_sb_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  assign LsuPlugin_logic_onAddress0_fromHp_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_3_ready;
  assign LsuPlugin_logic_onAddress0_arbiter_io_output_ready = (! execute_freeze_valid);
  assign execute_ctrl2_down_LsuL1_SEL_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  assign execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  always @(*) begin
    _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'bxxxxxxxx;
    case(LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size)
      2'b00 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h01;
      end
      2'b01 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h03;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'h0f;
      end
      default : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 8'hff;
      end
    endcase
  end

  assign execute_ctrl2_down_LsuL1_MASK_lane0 = (_zz_execute_ctrl2_down_LsuL1_MASK_lane0 <<< LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[2 : 0]);
  assign execute_ctrl2_down_LsuL1_SIZE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  assign execute_ctrl2_down_LsuL1_LOAD_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  assign execute_ctrl2_down_LsuL1_ATOMIC_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  assign execute_ctrl2_down_LsuL1_STORE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  assign execute_ctrl2_down_LsuL1_CLEAN_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  assign execute_ctrl2_down_LsuL1_INVALID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  assign execute_ctrl2_down_LsuL1_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign execute_ctrl2_down_LsuL1_FLUSH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_FLUSH);
  assign execute_ctrl2_down_Decode_STORE_ID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_ACCESS_1);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_STORE_BUFFER);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_LSU);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign execute_ctrl2_down_LsuPlugin_SB_PTR_lane0 = LsuPlugin_logic_storeBuffer_pop_payload_ptr;
  assign execute_ctrl2_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0 = LsuPlugin_logic_storeBuffer_pop_payload_op_data;
  assign execute_ctrl2_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0 = LsuPlugin_logic_storeBuffer_empty;
  assign execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign when_LsuPlugin_l546 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl3_up_LANE_SEL_lane0));
  assign when_LsuPlugin_l546_1 = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl4_up_LANE_SEL_lane0));
  assign execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = (|{((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b11) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 0] != 3'b000)),{((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b10) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0] != 2'b00)),((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b01) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[0 : 0] != 1'b0))}});
  assign execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = (((execute_ctrl3_down_AguPlugin_SEL_lane0 && execute_ctrl3_down_LsuL1_ATOMIC_lane0) && execute_ctrl3_down_LsuL1_STORE_lane0) && execute_ctrl3_down_LsuL1_LOAD_lane0);
  assign LsuPlugin_logic_onPma_cached_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_cached_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = LsuPlugin_logic_onPma_cached_rsp_fault;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = LsuPlugin_logic_onPma_cached_rsp_io;
  always @(*) begin
    execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = LsuPlugin_logic_onPma_io_rsp_fault;
    if(when_LsuPlugin_l569) begin
      execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = 1'b1;
    end
  end

  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = LsuPlugin_logic_onPma_io_rsp_io;
  assign when_LsuPlugin_l569 = (execute_ctrl3_down_LsuL1_ATOMIC_lane0 || execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0 = (((execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && (! execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault)) && (! execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0)) && (! execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onPma_addressExtension = 1'b0;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && 1'b0);
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = (execute_ctrl3_down_MMU_PAGE_FAULT_lane0 || (execute_ctrl3_down_AguPlugin_STORE_lane0 ? (! execute_ctrl3_down_MMU_ALLOW_WRITE_lane0) : (! execute_ctrl3_down_MMU_ALLOW_READ_lane0)));
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0 = ((((execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 || execute_ctrl3_down_MMU_ACCESS_FAULT_lane0) || execute_ctrl3_down_MMU_REFILL_lane0) || execute_ctrl3_down_MMU_HAZARD_lane0) || execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0);
  always @(*) begin
    LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(when_LsuPlugin_l759) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(when_LsuPlugin_l837) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_fenceTrap_valid) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
  end

  always @(*) begin
    LsuPlugin_logic_onCtrl_writeData = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuPlugin_logic_onCtrl_writeData[31 : 0] = execute_ctrl4_up_integer_RS2_lane0;
    if(execute_ctrl4_down_AguPlugin_FLOAT_lane0) begin
      LsuPlugin_logic_onCtrl_writeData[63 : 0] = execute_ctrl4_up_float_RS2_lane0;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) begin
      LsuPlugin_logic_onCtrl_writeData[31 : 0] = LsuPlugin_logic_onCtrl_rva_aluBuffer;
    end
  end

  assign when_LsuPlugin_l597 = (((((! LsuPlugin_logic_onCtrl_lsuTrap) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuPlugin_logic_onCtrl_io_doIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0);
  assign LsuPlugin_logic_bus_cmd_fire = (LsuPlugin_logic_bus_cmd_valid && LsuPlugin_logic_bus_cmd_ready);
  assign when_LsuPlugin_l601 = (! execute_freeze_valid);
  assign LsuPlugin_logic_bus_cmd_valid = (((LsuPlugin_logic_onCtrl_io_doItReg && (! LsuPlugin_logic_onCtrl_io_cmdSent)) && LsuPlugin_logic_onCtrl_io_allowIt) && (! LsuPlugin_logic_onCtrl_io_tooEarly));
  assign LsuPlugin_logic_bus_cmd_payload_write = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_size = execute_ctrl4_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_mask = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_io = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_fromHart = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_bus_rsp_toStream_valid = LsuPlugin_logic_bus_rsp_valid;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_error = LsuPlugin_logic_bus_rsp_payload_error;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_data = LsuPlugin_logic_bus_rsp_payload_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_fire = (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_ready);
  assign LsuPlugin_logic_bus_rsp_toStream_ready = (! LsuPlugin_logic_bus_rsp_toStream_rValid);
  assign LsuPlugin_logic_onCtrl_io_rsp_valid = LsuPlugin_logic_bus_rsp_toStream_rValid;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_error = LsuPlugin_logic_bus_rsp_toStream_rData_error;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_data = LsuPlugin_logic_bus_rsp_toStream_rData_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_ready = (! execute_freeze_valid);
  assign LsuPlugin_logic_onCtrl_io_freezeIt = (LsuPlugin_logic_onCtrl_io_doIt && (LsuPlugin_logic_onCtrl_io_tooEarly || ((! LsuPlugin_logic_onCtrl_io_rsp_valid) && LsuPlugin_logic_onCtrl_io_allowIt)));
  assign LsuPlugin_logic_onCtrl_loadData_input = (LsuPlugin_logic_onCtrl_io_cmdSent ? LsuPlugin_logic_onCtrl_io_rsp_payload_data : execute_ctrl4_down_LsuL1_READ_DATA_lane0);
  assign LsuPlugin_logic_onCtrl_loadData_splitted_0 = LsuPlugin_logic_onCtrl_loadData_input[7 : 0];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_1 = LsuPlugin_logic_onCtrl_loadData_input[15 : 8];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_2 = LsuPlugin_logic_onCtrl_loadData_input[23 : 16];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_3 = LsuPlugin_logic_onCtrl_loadData_input[31 : 24];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_4 = LsuPlugin_logic_onCtrl_loadData_input[39 : 32];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_5 = LsuPlugin_logic_onCtrl_loadData_input[47 : 40];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_6 = LsuPlugin_logic_onCtrl_loadData_input[55 : 48];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_7 = LsuPlugin_logic_onCtrl_loadData_input[63 : 56];
  always @(*) begin
    LsuPlugin_logic_onCtrl_loadData_shifted[7 : 0] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
    LsuPlugin_logic_onCtrl_loadData_shifted[15 : 8] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
    LsuPlugin_logic_onCtrl_loadData_shifted[23 : 16] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_4;
    LsuPlugin_logic_onCtrl_loadData_shifted[31 : 24] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_6;
    LsuPlugin_logic_onCtrl_loadData_shifted[39 : 32] = LsuPlugin_logic_onCtrl_loadData_splitted_4;
    LsuPlugin_logic_onCtrl_loadData_shifted[47 : 40] = LsuPlugin_logic_onCtrl_loadData_splitted_5;
    LsuPlugin_logic_onCtrl_loadData_shifted[55 : 48] = LsuPlugin_logic_onCtrl_loadData_splitted_6;
    LsuPlugin_logic_onCtrl_loadData_shifted[63 : 56] = LsuPlugin_logic_onCtrl_loadData_splitted_7;
  end

  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0 = LsuPlugin_logic_onCtrl_loadData_shifted;
  assign LsuPlugin_logic_onCtrl_storeData_mapping_0_1 = {8{LsuPlugin_logic_onCtrl_writeData[7 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_1_1 = {4{LsuPlugin_logic_onCtrl_writeData[15 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_2_1 = {2{LsuPlugin_logic_onCtrl_writeData[31 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_3_1 = {1{LsuPlugin_logic_onCtrl_writeData[63 : 0]}};
  always @(*) begin
    _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl4_down_LsuL1_SIZE_lane0)
      2'b00 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
      end
      2'b01 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
      end
      2'b10 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
      end
      default : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_3_1;
      end
    endcase
  end

  always @(*) begin
    execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
    if(execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0) begin
      execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = execute_ctrl4_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
    end
  end

  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0 = LsuPlugin_logic_onCtrl_scMiss;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_compare = execute_ctrl4_down_Decode_UOP_lane0[31 : 29];
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf = execute_ctrl4_down_Decode_UOP_lane0[27];
  assign LsuPlugin_logic_onCtrl_rva_alu_compare = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[2];
  assign LsuPlugin_logic_onCtrl_rva_alu_unsigned = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[1];
  assign LsuPlugin_logic_onCtrl_rva_alu_addSub = _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  assign LsuPlugin_logic_onCtrl_rva_alu_less = ((execute_ctrl4_down_integer_RS2_lane0[31] == LsuPlugin_logic_onCtrl_rva_srcBuffer[31]) ? LsuPlugin_logic_onCtrl_rva_alu_addSub[31] : (LsuPlugin_logic_onCtrl_rva_alu_unsigned ? LsuPlugin_logic_onCtrl_rva_srcBuffer[31] : execute_ctrl4_down_integer_RS2_lane0[31]));
  assign LsuPlugin_logic_onCtrl_rva_alu_selectRf = (_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf ? 1'b1 : (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare[0] ^ LsuPlugin_logic_onCtrl_rva_alu_less));
  assign switch_Misc_l245 = (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare | {_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf,2'b00});
  always @(*) begin
    case(switch_Misc_l245)
      3'b000 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = LsuPlugin_logic_onCtrl_rva_alu_addSub;
      end
      3'b001 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 ^ LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b010 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 | LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b011 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 & LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      default : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (LsuPlugin_logic_onCtrl_rva_alu_selectRf ? execute_ctrl4_down_integer_RS2_lane0 : LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
    endcase
  end

  assign LsuPlugin_logic_onCtrl_rva_alu_result = LsuPlugin_logic_onCtrl_rva_alu_raw;
  assign LsuPlugin_logic_onCtrl_rva_delay_0 = _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  assign LsuPlugin_logic_onCtrl_rva_delay_1 = _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  assign LsuPlugin_logic_onCtrl_rva_freezeIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) && (|{LsuPlugin_logic_onCtrl_rva_delay_1,LsuPlugin_logic_onCtrl_rva_delay_0}));
  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b0;
    if(when_LsuPlugin_l686) begin
      if(!execute_ctrl4_down_LsuL1_STORE_lane0) begin
        if(execute_ctrl4_down_LsuL1_ATOMIC_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b1;
        end
      end
    end
  end

  assign when_LsuPlugin_l686 = ((((((! execute_freeze_valid) && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && execute_ctrl4_down_LsuL1_SEL_lane0) && (! LsuPlugin_logic_onCtrl_lsuTrap)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign LsuPlugin_logic_onCtrl_scMiss = (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
  assign LsuL1_lockPort_valid = LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  assign LsuL1_lockPort_address = LsuPlugin_logic_onCtrl_rva_lrsc_address;
  assign when_LsuPlugin_l698 = ((! LsuPlugin_logic_onCtrl_rva_lrsc_age[5]) && (! execute_freeze_valid));
  assign when_LsuPlugin_l705 = (LsuPlugin_logic_onCtrl_rva_lrsc_age[5] || LsuPlugin_logic_onCtrl_io_cmdSent);
  assign when_LsuPlugin_l709 = (LsuPlugin_logic_onCtrl_rva_lrsc_capture && (LsuPlugin_logic_onCtrl_rva_lrsc_reserved || (6'h08 <= LsuPlugin_logic_onCtrl_rva_lrsc_age)));
  assign LsuPlugin_logic_onCtrl_wb_tag = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6];
  assign LsuPlugin_logic_onCtrl_wb_hits = {(LsuPlugin_logic_storeBuffer_slots_7_valid && (LsuPlugin_logic_storeBuffer_slots_7_tag == LsuPlugin_logic_onCtrl_wb_tag)),{(LsuPlugin_logic_storeBuffer_slots_6_valid && (LsuPlugin_logic_storeBuffer_slots_6_tag == LsuPlugin_logic_onCtrl_wb_tag)),{(LsuPlugin_logic_storeBuffer_slots_5_valid && (LsuPlugin_logic_storeBuffer_slots_5_tag == LsuPlugin_logic_onCtrl_wb_tag)),{(LsuPlugin_logic_storeBuffer_slots_4_valid && _zz_LsuPlugin_logic_onCtrl_wb_hits),{_zz_LsuPlugin_logic_onCtrl_wb_hits_1,{_zz_LsuPlugin_logic_onCtrl_wb_hits_2,_zz_LsuPlugin_logic_onCtrl_wb_hits_3}}}}}};
  assign LsuPlugin_logic_onCtrl_wb_hit = (|LsuPlugin_logic_onCtrl_wb_hits);
  assign LsuPlugin_logic_onCtrl_wb_compatibleOp = (((execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuL1_ATOMIC_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign LsuPlugin_logic_onCtrl_wb_notFull = ((! LsuPlugin_logic_storeBuffer_ops_full) && (LsuPlugin_logic_storeBuffer_slotsFree || LsuPlugin_logic_onCtrl_wb_hit));
  assign LsuPlugin_logic_onCtrl_wb_allowed = (LsuPlugin_logic_onCtrl_wb_notFull && LsuPlugin_logic_onCtrl_wb_compatibleOp);
  assign LsuPlugin_logic_onCtrl_wb_slotOh = (LsuPlugin_logic_onCtrl_wb_hits | ((! LsuPlugin_logic_onCtrl_wb_hit) ? LsuPlugin_logic_storeBuffer_slotsFreeFirst : 8'h0));
  assign LsuPlugin_logic_onCtrl_wb_loadHazard = (execute_ctrl4_down_LsuL1_LOAD_lane0 && LsuPlugin_logic_onCtrl_wb_hit);
  assign LsuPlugin_logic_onCtrl_wb_selfHazard = (execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0 && (execute_ctrl4_down_LsuPlugin_SB_PTR_lane0 != LsuPlugin_logic_storeBuffer_ops_freePtr));
  always @(*) begin
    LsuPlugin_logic_flushPort_valid = 1'b0;
    if(when_LsuPlugin_l865) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_flushPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_flushPort_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_flushPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane0;
  assign LsuPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    LsuPlugin_logic_trapPort_valid = 1'b0;
    if(when_LsuPlugin_l865) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_trapPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_trapPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane0;
  assign LsuPlugin_logic_trapPort_payload_tval = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  always @(*) begin
    LsuPlugin_logic_trapPort_payload_exception = 1'bx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(when_LsuPlugin_l759) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_fenceTrap_valid) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_code = 4'bxxxx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(when_LsuPlugin_l759) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b1101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
      if(when_LsuPlugin_l810) begin
        LsuPlugin_logic_trapPort_payload_code[3] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = {1'd0, _zz_LsuPlugin_logic_trapPort_payload_code};
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0011;
    end
    if(LsuPlugin_logic_onCtrl_fenceTrap_valid) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_arg = 2'b00;
    LsuPlugin_logic_trapPort_payload_arg[1 : 0] = (execute_ctrl4_down_LsuL1_STORE_lane0 ? 2'b01 : 2'b00);
  end

  assign LsuPlugin_logic_onCtrl_traps_accessFault = ((execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault ? (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_payload_error) : execute_ctrl4_down_LsuL1_FAULT_lane0) || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0);
  assign LsuPlugin_logic_onCtrl_traps_l1Failed = ((! execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault) && (execute_ctrl4_down_LsuL1_HAZARD_lane0 || ((execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && (execute_ctrl4_down_LsuL1_LOAD_lane0 || execute_ctrl4_down_LsuL1_STORE_lane0))));
  assign when_LsuPlugin_l759 = ((LsuPlugin_logic_onCtrl_traps_l1Failed || LsuPlugin_logic_onCtrl_wb_hit) && (! LsuPlugin_logic_onCtrl_wb_allowed));
  assign LsuPlugin_logic_onCtrl_traps_pmaFault = (execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault);
  assign when_LsuPlugin_l810 = (! execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0);
  always @(*) begin
    LsuPlugin_logic_storeBuffer_push_valid = 1'b0;
    if(when_LsuPlugin_l865) begin
      if(!LsuPlugin_logic_onCtrl_lsuTrap) begin
        if(when_LsuPlugin_l873) begin
          LsuPlugin_logic_storeBuffer_push_valid = 1'b1;
        end
      end
    end
  end

  assign LsuPlugin_logic_storeBuffer_push_payload_slotOh = LsuPlugin_logic_onCtrl_wb_slotOh;
  assign LsuPlugin_logic_storeBuffer_push_payload_tag = LsuPlugin_logic_onCtrl_wb_tag;
  assign LsuPlugin_logic_storeBuffer_push_payload_op_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuPlugin_logic_storeBuffer_push_payload_op_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign LsuPlugin_logic_storeBuffer_push_payload_op_size = execute_ctrl4_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_storeBuffer_push_payload_op_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign when_LsuPlugin_l837 = (execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign LsuPlugin_logic_onCtrl_fenceTrap_valid = ((execute_ctrl4_down_LsuL1_ATOMIC_lane0 || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0) && ((! LsuPlugin_logic_storeBuffer_empty) || (! execute_ctrl4_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0)));
  assign when_LsuPlugin_l865 = (execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0);
  assign when_LsuPlugin_l873 = (((LsuPlugin_logic_onCtrl_traps_l1Failed || LsuPlugin_logic_onCtrl_wb_hit) && LsuPlugin_logic_onCtrl_wb_allowed) && ((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)));
  assign when_LsuPlugin_l876 = (LsuPlugin_logic_onCtrl_wb_compatibleOp && (! LsuPlugin_logic_onCtrl_wb_notFull));
  assign LsuPlugin_logic_onCtrl_mmuNeeded = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign execute_ctrl4_down_LsuL1_ABORD_lane0 = (|{((LsuPlugin_logic_onCtrl_wb_loadHazard || ((! execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0) && LsuPlugin_logic_onCtrl_fenceTrap_valid)) || LsuPlugin_logic_onCtrl_wb_selfHazard),{(LsuPlugin_logic_onCtrl_mmuNeeded && execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0),{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (_zz_execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)),{(_zz_execute_ctrl4_down_LsuL1_ABORD_lane0_1 && execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault),{execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0,execute_ctrl4_down_LsuL1_HAZARD_lane0}}}}});
  assign execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0 = (|{(LsuPlugin_logic_onCtrl_wb_selfHazard || ((! execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0) && LsuPlugin_logic_onCtrl_wb_hit)),{((execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0)) && LsuPlugin_logic_onCtrl_scMiss),{execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0,{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0)),{execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0,{execute_ctrl4_down_LsuL1_FAULT_lane0,_zz_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0}}}}}});
  assign when_LsuPlugin_l905 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0) && ((execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 || execute_ctrl4_down_LsuL1_HAZARD_lane0) || execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0));
  assign when_LsuPlugin_l910 = (((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0) && (! execute_freeze_valid)) && (! LsuPlugin_logic_onCtrl_wb_selfHazard));
  assign when_LsuPlugin_l913 = (! execute_ctrl4_down_LsuL1_HAZARD_lane0);
  assign when_LsuPlugin_l263 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign when_LsuPlugin_l918 = (LsuPlugin_logic_storeBuffer_slots_0_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_1 = (LsuPlugin_logic_storeBuffer_slots_1_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_2 = (LsuPlugin_logic_storeBuffer_slots_2_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_3 = (LsuPlugin_logic_storeBuffer_slots_3_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_4 = (LsuPlugin_logic_storeBuffer_slots_4_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_5 = (LsuPlugin_logic_storeBuffer_slots_5_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_6 = (LsuPlugin_logic_storeBuffer_slots_6_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l918_7 = (LsuPlugin_logic_storeBuffer_slots_7_ptr == LsuPlugin_logic_storeBuffer_ops_freePtr);
  assign when_LsuPlugin_l259_1 = (|(LsuPlugin_logic_onCtrl_hartRegulation_refill & (~ LsuL1_REFILL_BUSY)));
  assign when_LsuPlugin_l949 = ((((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)) && execute_ctrl4_down_LsuL1_LOAD_lane0) && ((execute_ctrl4_down_LsuL1_HAZARD_lane0 || execute_ctrl4_down_LsuL1_MISS_lane0) || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0));
  assign when_LsuPlugin_l263_1 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign LsuPlugin_logic_onCtrl_commitProbeReq = ((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0);
  assign LsuPlugin_logic_commitProbe_valid = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (execute_ctrl4_down_AguPlugin_SEL_lane0 ? (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && ((! LsuPlugin_logic_onCtrl_lsuTrap) || (! LsuPlugin_logic_onCtrl_commitProbeToken))) : (execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 && execute_ctrl4_down_LsuL1_HAZARD_lane0)));
  assign LsuPlugin_logic_commitProbe_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  assign LsuPlugin_logic_commitProbe_payload_load = execute_ctrl4_down_LsuL1_LOAD_lane0;
  assign LsuPlugin_logic_commitProbe_payload_store = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_commitProbe_payload_trap = LsuPlugin_logic_onCtrl_lsuTrap;
  assign LsuPlugin_logic_commitProbe_payload_miss = ((execute_ctrl4_down_LsuL1_MISS_lane0 && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0));
  assign LsuPlugin_logic_commitProbe_payload_io = execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  assign LsuPlugin_logic_commitProbe_payload_prefetchFailed = execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign LsuPlugin_logic_commitProbe_payload_pc = execute_ctrl4_down_PC_lane0;
  assign LsuPlugin_logic_iwb_valid = (execute_ctrl4_down_AguPlugin_SEL_lane0 && (! execute_ctrl4_down_AguPlugin_FLOAT_lane0));
  always @(*) begin
    LsuPlugin_logic_iwb_payload = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0[31:0];
    if(when_LsuPlugin_l974) begin
      LsuPlugin_logic_iwb_payload[0] = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
      LsuPlugin_logic_iwb_payload[7 : 1] = 7'h0;
    end
  end

  assign when_LsuPlugin_l974 = (execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0));
  assign LsuPlugin_logic_fpwb_valid = (execute_ctrl4_down_AguPlugin_SEL_lane0 && execute_ctrl4_down_AguPlugin_FLOAT_lane0);
  always @(*) begin
    LsuPlugin_logic_fpwb_payload = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    if(when_LsuPlugin_l982) begin
      LsuPlugin_logic_fpwb_payload[63 : 32] = 32'hffffffff;
    end
  end

  assign when_LsuPlugin_l982 = (execute_ctrl4_down_AguPlugin_SIZE_lane0 == 2'b10);
  assign LsuPlugin_logic_onWb_storeFire = ((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onWb_storeBroadcast = (((((((execute_ctrl4_down_isReady && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuL1_ABORD_lane0)) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)) && (! execute_ctrl4_down_LsuL1_HAZARD_lane0));
  always @(*) begin
    LsuPlugin_logic_storeBuffer_ops_pip_node_0_ready = LsuPlugin_logic_storeBuffer_ops_pip_node_1_ready;
    if(when_StageLink_l71_1) begin
      LsuPlugin_logic_storeBuffer_ops_pip_node_0_ready = 1'b1;
    end
  end

  assign when_StageLink_l71_1 = (! LsuPlugin_logic_storeBuffer_ops_pip_node_1_isValid);
  always @(*) begin
    LsuPlugin_logic_storeBuffer_ops_pip_node_1_ready = LsuPlugin_logic_storeBuffer_ops_pip_node_2_ready;
    if(when_StageLink_l71_2) begin
      LsuPlugin_logic_storeBuffer_ops_pip_node_1_ready = 1'b1;
    end
  end

  assign when_StageLink_l71_2 = (! LsuPlugin_logic_storeBuffer_ops_pip_node_2_isValid);
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_0_isFiring = (LsuPlugin_logic_storeBuffer_ops_pip_node_0_isValid && LsuPlugin_logic_storeBuffer_ops_pip_node_0_isReady);
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_0_isValid = LsuPlugin_logic_storeBuffer_ops_pip_node_0_valid;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_0_isReady = LsuPlugin_logic_storeBuffer_ops_pip_node_0_ready;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_isValid = LsuPlugin_logic_storeBuffer_ops_pip_node_1_valid;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_1_isReady = LsuPlugin_logic_storeBuffer_ops_pip_node_1_ready;
  assign LsuPlugin_logic_storeBuffer_ops_pip_node_2_isValid = LsuPlugin_logic_storeBuffer_ops_pip_node_2_valid;
  assign FpuPackerPlugin_logic_s0_remapped_0_mode = FpuUnpackerPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_0_quiet = FpuUnpackerPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_0_sign = FpuUnpackerPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_0_exponent = {7'd0, FpuUnpackerPlugin_logic_packPort_cmd_value_exponent};
  assign FpuPackerPlugin_logic_s0_remapped_0_mantissa = FpuUnpackerPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuPackerPlugin_logic_s0_remapped_1_mode = FpuMulPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_1_quiet = FpuMulPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_1_sign = FpuMulPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_1_exponent = _zz_FpuPackerPlugin_logic_s0_remapped_1_exponent;
  assign FpuPackerPlugin_logic_s0_remapped_1_mantissa = FpuMulPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuPackerPlugin_logic_s0_remapped_2_mode = FpuSqrtPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_2_quiet = FpuSqrtPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_2_sign = FpuSqrtPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_2_exponent = _zz_FpuPackerPlugin_logic_s0_remapped_2_exponent;
  assign FpuPackerPlugin_logic_s0_remapped_2_mantissa = FpuSqrtPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuPackerPlugin_logic_s0_remapped_3_mode = FpuXxPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_3_quiet = FpuXxPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_3_sign = FpuXxPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_3_exponent = _zz_FpuPackerPlugin_logic_s0_remapped_3_exponent;
  assign FpuPackerPlugin_logic_s0_remapped_3_mantissa = FpuXxPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuPackerPlugin_logic_s0_remapped_4_mode = FpuDivPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_4_quiet = FpuDivPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_4_sign = FpuDivPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_4_exponent = _zz_FpuPackerPlugin_logic_s0_remapped_4_exponent;
  assign FpuPackerPlugin_logic_s0_remapped_4_mantissa = FpuDivPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuPackerPlugin_logic_s0_remapped_5_mode = FpuAddSharedPlugin_logic_packPort_cmd_value_mode;
  assign FpuPackerPlugin_logic_s0_remapped_5_quiet = FpuAddSharedPlugin_logic_packPort_cmd_value_quiet;
  assign FpuPackerPlugin_logic_s0_remapped_5_sign = FpuAddSharedPlugin_logic_packPort_cmd_value_sign;
  assign FpuPackerPlugin_logic_s0_remapped_5_exponent = _zz_FpuPackerPlugin_logic_s0_remapped_5_exponent;
  assign FpuPackerPlugin_logic_s0_remapped_5_mantissa = FpuAddSharedPlugin_logic_packPort_cmd_value_mantissa;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid = (|FpuUnpackerPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid_1 = (|FpuMulPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid_2 = (|FpuSqrtPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid_3 = (|FpuXxPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid_4 = (|FpuDivPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_valid_5 = (|FpuAddSharedPlugin_logic_packPort_cmd_at);
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet = {_zz_FpuPackerPlugin_logic_pip_node_0_valid_5,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_4,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_3,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_2,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_1,_zz_FpuPackerPlugin_logic_pip_node_0_valid}}}}};
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1 = ((((_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_1 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_4) | (_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_5 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_6 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_9)) | ((_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_10 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_11 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_14) | (_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_15 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_16 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_19))) | ((_zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[4] ? {FpuPackerPlugin_logic_s0_remapped_4_mantissa,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_20} : 71'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet[5] ? {FpuPackerPlugin_logic_s0_remapped_5_mantissa,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1_23} : 71'h0)));
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1 = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1[1 : 0];
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode_1;
  assign FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode;
  assign FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1[2];
  assign FpuPackerPlugin_logic_pip_node_0_s0_VALUE_sign = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet_1[3];
  assign FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_exponent;
  assign FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa = _zz_FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa[53 : 0];
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1 = ((((_zz_FpuPackerPlugin_logic_pip_node_0_valid ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_1) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_1 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_2 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_3)) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_2 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_4 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_5) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_3 ? _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_6 : _zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1_7))) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_4 ? FpuDivPlugin_logic_packPort_cmd_format : 1'b0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_5 ? FpuAddSharedPlugin_logic_packPort_cmd_format : 1'b0)));
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT_1;
  assign FpuPackerPlugin_logic_pip_node_0_s0_FORMAT = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FORMAT;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1 = ((((_zz_FpuPackerPlugin_logic_pip_node_0_valid ? FpuUnpackerPlugin_logic_packPort_cmd_roundMode : 3'b000) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_1 ? FpuMulPlugin_logic_packPort_cmd_roundMode : 3'b000)) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_2 ? FpuSqrtPlugin_logic_packPort_cmd_roundMode : 3'b000) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_3 ? FpuXxPlugin_logic_packPort_cmd_roundMode : 3'b000))) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_4 ? FpuDivPlugin_logic_packPort_cmd_roundMode : 3'b000) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_5 ? FpuAddSharedPlugin_logic_packPort_cmd_roundMode : 3'b000)));
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE = _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE_1;
  assign FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE = _zz_FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE;
  assign _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX = ((((_zz_FpuPackerPlugin_logic_pip_node_0_valid ? {_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_1} : 5'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_1 ? {_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_4,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_5} : 5'h0)) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_2 ? {_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_8,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_9} : 5'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_3 ? {_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_12,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_13} : 5'h0))) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_4 ? {FpuDivPlugin_logic_packPort_cmd_flags_NV,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_16,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_17}} : 5'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_5 ? {FpuAddSharedPlugin_logic_packPort_cmd_flags_NV,{_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_20,_zz__zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX_21}} : 5'h0)));
  assign FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX[0];
  assign FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_UF = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX[1];
  assign FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_OF = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX[2];
  assign FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_DZ = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX[3];
  assign FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NV = _zz_FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX[4];
  assign FpuPackerPlugin_logic_pip_node_0_Decode_UOP_ID = ((((_zz_FpuPackerPlugin_logic_pip_node_0_valid ? FpuUnpackerPlugin_logic_packPort_cmd_uopId : 16'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_1 ? FpuMulPlugin_logic_packPort_cmd_uopId : 16'h0)) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_2 ? FpuSqrtPlugin_logic_packPort_cmd_uopId : 16'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_3 ? FpuXxPlugin_logic_packPort_cmd_uopId : 16'h0))) | ((_zz_FpuPackerPlugin_logic_pip_node_0_valid_4 ? FpuDivPlugin_logic_packPort_cmd_uopId : 16'h0) | (_zz_FpuPackerPlugin_logic_pip_node_0_valid_5 ? FpuAddSharedPlugin_logic_packPort_cmd_uopId : 16'h0)));
  assign FpuPackerPlugin_logic_pip_node_0_valid = (|{_zz_FpuPackerPlugin_logic_pip_node_0_valid_5,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_4,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_3,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_2,{_zz_FpuPackerPlugin_logic_pip_node_0_valid_1,_zz_FpuPackerPlugin_logic_pip_node_0_valid}}}}});
  assign _zz_49 = 3'b000;
  assign _zz_50 = 3'b001;
  assign _zz_51 = 3'b001;
  assign _zz_52 = 3'b010;
  assign _zz_53 = 3'b001;
  assign _zz_54 = 3'b010;
  assign _zz_55 = 3'b010;
  assign _zz_56 = 3'b011;
  always @(*) begin
    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[0] = (|{FpuDivPlugin_logic_packPort_cmd_at[0],{FpuSqrtPlugin_logic_packPort_cmd_at[0],FpuUnpackerPlugin_logic_packPort_cmd_at[0]}});
    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[1] = (|FpuMulPlugin_logic_packPort_cmd_at[0]);
    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[2] = (|FpuXxPlugin_logic_packPort_cmd_at[0]);
    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[3] = (|FpuAddSharedPlugin_logic_packPort_cmd_at[0]);
    FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH[4] = (|FpuAddSharedPlugin_logic_packPort_cmd_at[1]);
  end

  assign FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL = _zz_FpuPackerPlugin_logic_pip_node_0_s0_EXP_SUBNORMAL;
  assign FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE = (($signed(_zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE) <= $signed(_zz_FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE_1)) && (FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode == FloatMode_NORMAL));
  always @(*) begin
    FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED = FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mantissa;
    if(FpuPackerPlugin_logic_pip_node_1_s0_subnormal_ENABLE) begin
      FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED = FpuPackerPlugin_logic_s1_subnormal_manShifter;
    end
  end

  assign _zz_when_AFix_l1168_1 = _zz__zz_when_AFix_l1168_1_1;
  assign when_AFix_l1168_1 = _zz_when_AFix_l1168_1[12];
  always @(*) begin
    if(when_AFix_l1168_1) begin
      _zz_FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE = 13'h0;
    end else begin
      _zz_FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE = _zz_when_AFix_l1168_1;
    end
  end

  assign FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE = (_zz_FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE + 13'h0001);
  assign when_UInt_l119_1 = (|FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE[12 : 6]);
  always @(*) begin
    if(when_UInt_l119_1) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShift = 6'h3f;
    end else begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShift = FpuPackerPlugin_logic_pip_node_1_s1_subnormal_EXP_DIF_PLUS_ONE[5 : 0];
    end
  end

  assign _zz_when_Utils_l1585_15 = {1'b1,FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mantissa};
  always @(*) begin
    _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b0;
    if(when_Utils_l1585_7) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
    if(when_Utils_l1585_8) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
    if(when_Utils_l1585_9) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
    if(when_Utils_l1585_10) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
    if(when_Utils_l1585_11) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
    if(when_Utils_l1585_12) begin
      _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_1 = 1'b1;
    end
  end

  assign when_Utils_l1585_7 = (FpuPackerPlugin_logic_s1_subnormal_manShift[0] && (_zz_when_Utils_l1585_15[0 : 0] != 1'b0));
  assign when_Utils_l1585_8 = (FpuPackerPlugin_logic_s1_subnormal_manShift[1] && (_zz_when_Utils_l1585_7[1 : 0] != 2'b00));
  assign when_Utils_l1585_9 = (FpuPackerPlugin_logic_s1_subnormal_manShift[2] && (_zz_when_Utils_l1585_6[3 : 0] != 4'b0000));
  assign when_Utils_l1585_10 = (FpuPackerPlugin_logic_s1_subnormal_manShift[3] && (_zz_when_Utils_l1585_5[7 : 0] != 8'h0));
  assign when_Utils_l1585_11 = (FpuPackerPlugin_logic_s1_subnormal_manShift[4] && (_zz_when_Utils_l1585_4[15 : 0] != 16'h0));
  assign when_Utils_l1585_12 = (FpuPackerPlugin_logic_s1_subnormal_manShift[5] && (_zz_when_Utils_l1585_3[31 : 0] != 32'h0));
  assign FpuPackerPlugin_logic_s1_subnormal_freezeIt = ((FpuPackerPlugin_logic_pip_node_1_isValid && FpuPackerPlugin_logic_pip_node_1_s0_subnormal_ENABLE) && (FpuPackerPlugin_logic_s1_subnormal_counter != 2'b10));
  assign when_FpuPackerPlugin_l134 = (! execute_freeze_valid);
  assign FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted = ((FpuPackerPlugin_logic_pip_node_1_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED[1 : 0] : (FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED[30 : 29] | _zz_FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted));
  assign FpuPackerPlugin_logic_pip_node_1_s1_manLsb = ((FpuPackerPlugin_logic_pip_node_1_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED[2] : FpuPackerPlugin_logic_pip_node_1_s1_MAN_SHIFTED[31]);
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE)
      FpuRoundMode_RNE : begin
        _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = (FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted[1] && (FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted[0] || FpuPackerPlugin_logic_pip_node_1_s1_manLsb));
      end
      FpuRoundMode_RTZ : begin
        _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = 1'b0;
      end
      FpuRoundMode_RDN : begin
        _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = ((FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted != 2'b00) && FpuPackerPlugin_logic_pip_node_1_s0_VALUE_sign);
      end
      FpuRoundMode_RUP : begin
        _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = ((FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted != 2'b00) && (! FpuPackerPlugin_logic_pip_node_1_s0_VALUE_sign));
      end
      default : begin
        _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted[1];
      end
    endcase
  end

  assign FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR = ((FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode == FloatMode_NORMAL) && _zz_FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR);
  assign FpuPackerPlugin_logic_s1_incrBy = ((FpuPackerPlugin_logic_pip_node_1_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? 30'h00000001 : _zz_FpuPackerPlugin_logic_s1_incrBy);
  assign FpuPackerPlugin_logic_s1_manIncrWithCarry = ({1'b0,_zz_FpuPackerPlugin_logic_s1_manIncrWithCarry} + _zz_FpuPackerPlugin_logic_s1_manIncrWithCarry_1);
  assign FpuPackerPlugin_logic_s1_MAN_CARRY = FpuPackerPlugin_logic_s1_manIncrWithCarry[52];
  assign FpuPackerPlugin_logic_s1_MAN_INCR = FpuPackerPlugin_logic_s1_manIncrWithCarry[51 : 0];
  assign FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR = _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_INCR;
  assign FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT = _zz_FpuPackerPlugin_logic_pip_node_1_s1_EXP_RESULT;
  assign FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT = (FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR ? FpuPackerPlugin_logic_s1_MAN_INCR : _zz_FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT);
  assign FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL = (! _zz_FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL[12]);
  assign FpuPackerPlugin_logic_pip_node_2_s2_EXP = _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP;
  assign FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX = _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MAX;
  assign FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN = _zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_MIN;
  assign FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW = ($signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) < $signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW_2));
  assign FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW = ($signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) < $signed(_zz_FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW_1));
  assign FpuPackerPlugin_logic_s2_tinyRound = ((FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? {FpuPackerPlugin_logic_s2_mr[1],(|FpuPackerPlugin_logic_s2_mr[0 : 0])} : {FpuPackerPlugin_logic_s2_mr[30],(|FpuPackerPlugin_logic_s2_mr[29 : 0])});
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE)
      FpuRoundMode_RNE : begin
        _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr = (FpuPackerPlugin_logic_s2_tinyRound[1] && (FpuPackerPlugin_logic_s2_tinyRound[0] || FpuPackerPlugin_logic_pip_node_2_s1_manLsb));
      end
      FpuRoundMode_RTZ : begin
        _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr = 1'b0;
      end
      FpuRoundMode_RDN : begin
        _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr = ((FpuPackerPlugin_logic_s2_tinyRound != 2'b00) && FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign);
      end
      FpuRoundMode_RUP : begin
        _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr = ((FpuPackerPlugin_logic_s2_tinyRound != 2'b00) && (! FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign));
      end
      default : begin
        _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr = FpuPackerPlugin_logic_s2_tinyRound[1];
      end
    endcase
  end

  assign FpuPackerPlugin_logic_s2_tinyRoundingIncr = ((FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode == FloatMode_NORMAL) && _zz_FpuPackerPlugin_logic_s2_tinyRoundingIncr);
  assign FpuPackerPlugin_logic_s2_tinyOverflow = (((FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1) ? (&FpuPackerPlugin_logic_s2_mr[53 : 2]) : (&FpuPackerPlugin_logic_s2_mr[53 : 31])) && FpuPackerPlugin_logic_s2_tinyRoundingIncr);
  always @(*) begin
    FpuPackerPlugin_logic_s2_expSet = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
        FpuPackerPlugin_logic_s2_expSet = 1'b1;
      end
      FloatMode_NAN : begin
        FpuPackerPlugin_logic_s2_expSet = 1'b1;
      end
      default : begin
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(!when_FpuPackerPlugin_l224) begin
            FpuPackerPlugin_logic_s2_expSet = 1'b1;
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_expZero = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
        FpuPackerPlugin_logic_s2_expZero = 1'b1;
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(!FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) begin
            if(when_FpuPackerPlugin_l241) begin
              FpuPackerPlugin_logic_s2_expZero = 1'b1;
            end else begin
              FpuPackerPlugin_logic_s2_expZero = 1'b1;
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_expMax = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(when_FpuPackerPlugin_l224) begin
            FpuPackerPlugin_logic_s2_expMax = 1'b1;
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_manZero = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
        FpuPackerPlugin_logic_s2_manZero = 1'b1;
      end
      FloatMode_INF : begin
        FpuPackerPlugin_logic_s2_manZero = 1'b1;
      end
      FloatMode_NAN : begin
        FpuPackerPlugin_logic_s2_manZero = 1'b1;
      end
      default : begin
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(!when_FpuPackerPlugin_l224) begin
            FpuPackerPlugin_logic_s2_manZero = 1'b1;
          end
        end else begin
          if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) begin
            if(!when_FpuPackerPlugin_l241) begin
              FpuPackerPlugin_logic_s2_manZero = 1'b1;
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_manSet = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(when_FpuPackerPlugin_l224) begin
            FpuPackerPlugin_logic_s2_manSet = 1'b1;
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_manOne = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(!FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) begin
            if(when_FpuPackerPlugin_l241) begin
              FpuPackerPlugin_logic_s2_manOne = 1'b1;
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_manQuiet = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
        FpuPackerPlugin_logic_s2_manQuiet = FpuPackerPlugin_logic_pip_node_2_s0_VALUE_quiet;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_positive = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
        FpuPackerPlugin_logic_s2_positive = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_nx = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(when_FpuPackerPlugin_l208) begin
          FpuPackerPlugin_logic_s2_nx = 1'b1;
        end
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          FpuPackerPlugin_logic_s2_nx = 1'b1;
        end else begin
          if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) begin
            FpuPackerPlugin_logic_s2_nx = 1'b1;
          end
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_of = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          FpuPackerPlugin_logic_s2_of = 1'b1;
        end
      end
    endcase
  end

  always @(*) begin
    FpuPackerPlugin_logic_s2_uf = 1'b0;
    case(FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode)
      FloatMode_ZERO : begin
      end
      FloatMode_INF : begin
      end
      FloatMode_NAN : begin
      end
      default : begin
        if(when_FpuPackerPlugin_l208) begin
          if(when_FpuPackerPlugin_l210) begin
            FpuPackerPlugin_logic_s2_uf = 1'b1;
          end
        end
        if(!FpuPackerPlugin_logic_pip_node_2_s2_EXP_OVERFLOW) begin
          if(FpuPackerPlugin_logic_pip_node_2_s2_EXP_UNDERFLOW) begin
            FpuPackerPlugin_logic_s2_uf = 1'b1;
          end
        end
      end
    endcase
  end

  assign when_FpuPackerPlugin_l208 = (FpuPackerPlugin_logic_pip_node_2_s1_roundAdjusted != 2'b00);
  assign when_FpuPackerPlugin_l210 = (FpuPackerPlugin_logic_pip_node_2_s2_SUBNORMAL_FINAL || (FpuPackerPlugin_logic_pip_node_2_s0_subnormal_ENABLE && (! FpuPackerPlugin_logic_s2_tinyOverflow)));
  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE)
      FpuRoundMode_RNE : begin
        when_FpuPackerPlugin_l224 = 1'b0;
      end
      FpuRoundMode_RTZ : begin
        when_FpuPackerPlugin_l224 = 1'b1;
      end
      FpuRoundMode_RDN : begin
        when_FpuPackerPlugin_l224 = (! FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign);
      end
      FpuRoundMode_RUP : begin
        when_FpuPackerPlugin_l224 = FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign;
      end
      default : begin
        when_FpuPackerPlugin_l224 = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE)
      FpuRoundMode_RNE : begin
        _zz_when_FpuPackerPlugin_l241 = 1'b0;
      end
      FpuRoundMode_RTZ : begin
        _zz_when_FpuPackerPlugin_l241 = 1'b0;
      end
      FpuRoundMode_RDN : begin
        _zz_when_FpuPackerPlugin_l241 = FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign;
      end
      FpuRoundMode_RUP : begin
        _zz_when_FpuPackerPlugin_l241 = (! FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign);
      end
      default : begin
        _zz_when_FpuPackerPlugin_l241 = 1'b0;
      end
    endcase
  end

  assign when_FpuPackerPlugin_l241 = (_zz_when_FpuPackerPlugin_l241 || FpuPackerPlugin_logic_pip_node_2_s1_ROUNDING_INCR);
  assign FpuPackerPlugin_wb_at_2_valid = FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH[0];
  assign FpuPackerPlugin_wb_at_2_payload = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_wb_at_5_valid = FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH[1];
  assign FpuPackerPlugin_wb_at_5_payload = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_wb_at_3_valid = FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH[2];
  assign FpuPackerPlugin_wb_at_3_payload = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_wb_at_6_valid = FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH[3];
  assign FpuPackerPlugin_wb_at_6_payload = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_wb_at_9_valid = FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH[4];
  assign FpuPackerPlugin_wb_at_9_payload = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_logic_s2_fpWriter_valid = ((|FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH) && FpuPackerPlugin_logic_pip_node_2_valid);
  assign FpuPackerPlugin_logic_s2_fpWriter_payload_data = FpuPackerPlugin_logic_s2_fwb_value;
  assign FpuPackerPlugin_logic_s2_fpWriter_payload_uopId = FpuPackerPlugin_logic_pip_node_2_Decode_UOP_ID;
  assign FpuPackerPlugin_logic_flagsWb_ats = (FpuPackerPlugin_logic_pip_node_2_valid ? FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH : 5'h0);
  assign FpuPackerPlugin_logic_flagsWb_flags_NX = (FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NX || FpuPackerPlugin_logic_s2_nx);
  assign FpuPackerPlugin_logic_flagsWb_flags_UF = (FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_UF || FpuPackerPlugin_logic_s2_uf);
  assign FpuPackerPlugin_logic_flagsWb_flags_OF = (FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_OF || FpuPackerPlugin_logic_s2_of);
  assign FpuPackerPlugin_logic_flagsWb_flags_DZ = FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_DZ;
  assign FpuPackerPlugin_logic_flagsWb_flags_NV = FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NV;
  assign when_Misc_l22 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  always @(*) begin
    if(when_Misc_l22) begin
      FpuPackerPlugin_logic_s2_fwb_value = {{FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign,_zz_FpuPackerPlugin_logic_s2_fwb_value},FpuPackerPlugin_logic_pip_node_2_s1_MAN_RESULT};
    end else begin
      FpuPackerPlugin_logic_s2_fwb_value[31 : 0] = {{FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign,FpuPackerPlugin_logic_pip_node_2_s2_EXP[7 : 0]},FpuPackerPlugin_logic_pip_node_2_s1_MAN_RESULT[51 : 29]};
      FpuPackerPlugin_logic_s2_fwb_value[63 : 32] = 32'hffffffff;
    end
    if(FpuPackerPlugin_logic_s2_expZero) begin
      if(when_Misc_l22_1) begin
        FpuPackerPlugin_logic_s2_fwb_value[62 : 52] = 11'h0;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[30 : 23] = 8'h0;
      end
    end
    if(FpuPackerPlugin_logic_s2_expSet) begin
      if(when_Misc_l22_2) begin
        FpuPackerPlugin_logic_s2_fwb_value[62 : 52] = 11'h7ff;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[30 : 23] = 8'hff;
      end
    end
    if(FpuPackerPlugin_logic_s2_expMax) begin
      if(when_Misc_l22_3) begin
        FpuPackerPlugin_logic_s2_fwb_value[62 : 52] = 11'h7fe;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[30 : 23] = 8'hfe;
      end
    end
    if(FpuPackerPlugin_logic_s2_manZero) begin
      if(when_Misc_l22_4) begin
        FpuPackerPlugin_logic_s2_fwb_value[51 : 0] = 52'h0;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[22 : 0] = 23'h0;
      end
    end
    if(FpuPackerPlugin_logic_s2_manOne) begin
      if(when_Misc_l22_5) begin
        FpuPackerPlugin_logic_s2_fwb_value[51 : 0] = 52'h0000000000001;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[22 : 0] = 23'h000001;
      end
    end
    if(FpuPackerPlugin_logic_s2_manSet) begin
      if(when_Misc_l22_6) begin
        FpuPackerPlugin_logic_s2_fwb_value[51 : 0] = 52'hfffffffffffff;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[22 : 0] = 23'h7fffff;
      end
    end
    if(FpuPackerPlugin_logic_s2_manQuiet) begin
      if(when_Misc_l22_7) begin
        FpuPackerPlugin_logic_s2_fwb_value[51] = 1'b1;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[22] = 1'b1;
      end
    end
    if(FpuPackerPlugin_logic_s2_positive) begin
      if(when_Misc_l22_8) begin
        FpuPackerPlugin_logic_s2_fwb_value[63] = 1'b0;
      end else begin
        FpuPackerPlugin_logic_s2_fwb_value[31] = 1'b0;
      end
    end
    if(when_FpuPackerPlugin_l309) begin
      FpuPackerPlugin_logic_s2_fwb_value[63 : 32] = 32'hffffffff;
    end
  end

  assign when_Misc_l22_1 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_2 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_3 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_4 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_5 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_6 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_7 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_8 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_FpuPackerPlugin_l309 = (FpuPackerPlugin_logic_pip_node_2_s0_FORMAT == FpuFormat_FpuCmpPlugin_logic_f32_1);
  assign FpuPackerPlugin_logic_pip_node_2_ready = (! execute_freeze_valid);
  assign FpuPackerPlugin_logic_pip_node_0_ready = FpuPackerPlugin_logic_pip_node_1_ready;
  assign FpuPackerPlugin_logic_pip_node_1_ready = FpuPackerPlugin_logic_pip_node_2_ready;
  assign FpuPackerPlugin_logic_pip_node_0_isValid = FpuPackerPlugin_logic_pip_node_0_valid;
  assign FpuPackerPlugin_logic_pip_node_0_isReady = FpuPackerPlugin_logic_pip_node_0_ready;
  assign FpuPackerPlugin_logic_pip_node_1_isValid = FpuPackerPlugin_logic_pip_node_1_valid;
  assign FpuPackerPlugin_logic_pip_node_1_isReady = FpuPackerPlugin_logic_pip_node_1_ready;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) == $signed(execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0));
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 != execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign early0_BranchPlugin_logic_alu_expectedMsb = 1'b0;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l245_1 = execute_ctrl2_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l245_1)
      3'b000 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl2_down_early0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 ? execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 != execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_needFix = ((early0_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 && execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_BranchPlugin_SEL_lane0) && early0_BranchPlugin_logic_jumpLogic_needFix);
  assign early0_BranchPlugin_logic_jumpLogic_history_slice = execute_ctrl2_down_PC_lane0[2 : 1];
  assign early0_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l213 = ((early0_BranchPlugin_logic_jumpLogic_history_slice < 2'b00) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[0]);
  assign when_BranchPlugin_l213_1 = ((early0_BranchPlugin_logic_jumpLogic_history_slice < 2'b01) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[1]);
  assign when_BranchPlugin_l213_2 = ((early0_BranchPlugin_logic_jumpLogic_history_slice < 2'b10) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[2]);
  assign when_BranchPlugin_l218 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_history_next = early0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  assign early0_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  assign early0_BranchPlugin_logic_pcPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_historyPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_historyPort_payload_history = early0_BranchPlugin_logic_jumpLogic_history_next;
  assign early0_BranchPlugin_logic_historyPort_payload_age = execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_flushPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0 : 0] != 1'b0) && execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early0_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl2_down_Decode_UOP_lane0[11 : 7] == execute_ctrl2_down_Decode_UOP_lane0[19 : 15]);
  assign early0_BranchPlugin_logic_wb_valid = execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  assign early0_BranchPlugin_logic_wb_payload = execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1 = ($signed(execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1) == $signed(execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1));
  assign execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1 != execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1);
  assign early1_BranchPlugin_logic_alu_expectedMsb = 1'b0;
  assign execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1 = ((execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l245_2 = execute_ctrl2_down_Decode_UOP_lane1[14 : 12];
  always @(*) begin
    casez(switch_Misc_l245_2)
      3'b000 : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1;
      end
      3'b001 : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1);
      end
      3'b1?1 : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! execute_ctrl2_down_early1_SrcPlugin_LESS_lane1);
      end
      default : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
      end
    endcase
  end

  assign execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = _zz_execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  assign execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1 = (execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 ? execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 : execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1 != execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_needFix = ((early1_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 && execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1)) || execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl2_up_LANE_SEL_lane1 && execute_ctrl2_down_early1_BranchPlugin_SEL_lane1) && early1_BranchPlugin_logic_jumpLogic_needFix);
  assign early1_BranchPlugin_logic_jumpLogic_history_slice = execute_ctrl2_down_PC_lane1[2 : 1];
  assign early1_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
  assign when_BranchPlugin_l213_3 = ((early1_BranchPlugin_logic_jumpLogic_history_slice < 2'b00) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[0]);
  assign when_BranchPlugin_l213_4 = ((early1_BranchPlugin_logic_jumpLogic_history_slice < 2'b01) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[1]);
  assign when_BranchPlugin_l213_5 = ((early1_BranchPlugin_logic_jumpLogic_history_slice < 2'b10) && execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[2]);
  assign when_BranchPlugin_l218_1 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign early1_BranchPlugin_logic_jumpLogic_history_next = early1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  assign early1_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
  assign early1_BranchPlugin_logic_pcPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  assign early1_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  assign early1_BranchPlugin_logic_pcPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_historyPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_historyPort_payload_history = early1_BranchPlugin_logic_jumpLogic_history_next;
  assign early1_BranchPlugin_logic_historyPort_payload_age = execute_ctrl2_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_flushPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign early1_BranchPlugin_logic_flushPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1 = ((execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0 : 0] != 1'b0) && execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl2_down_early1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 = (execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early1_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl2_down_Decode_UOP_lane1[11 : 7] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane1[11 : 7] == 5'h01)});
  assign early1_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl2_down_Decode_UOP_lane1[19 : 15] == 5'h05),(execute_ctrl2_down_Decode_UOP_lane1[19 : 15] == 5'h01)});
  assign early1_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl2_down_Decode_UOP_lane1[11 : 7] == execute_ctrl2_down_Decode_UOP_lane1[19 : 15]);
  assign early1_BranchPlugin_logic_wb_valid = execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
  assign early1_BranchPlugin_logic_wb_payload = execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign PmpPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign PmpPlugin_logic_instructionShouldHit = (! PmpPlugin_logic_isMachine);
  assign PmpPlugin_logic_dataShouldHit = ((! PmpPlugin_logic_isMachine) || (PrivilegedPlugin_logic_harts_0_m_status_mprv && (PrivilegedPlugin_logic_harts_0_m_status_mpp != 2'b11)));
  assign FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || 1'b0);
  assign FetchL1Plugin_logic_pmpPort_logic_torCmpAddress = (fetch_logic_ctrls_1_down_MMU_TRANSLATED >>> 4'd12);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT = ((PmpPlugin_logic_instructionShouldHit && 1'b1) || (FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort && (1'b0 || 1'b0)));
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT = 1'b0;
  assign LsuPlugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign LsuPlugin_logic_pmpPort_logic_torCmpAddress = (execute_ctrl3_down_MMU_TRANSLATED_lane0 >>> 4'd12);
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 = ((PmpPlugin_logic_instructionShouldHit && 1'b0) || (LsuPlugin_logic_pmpPort_logic_dataShouldHitPort && (execute_ctrl2_down_LsuL1_LOAD_lane0 || execute_ctrl2_down_LsuL1_STORE_lane0)));
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 = 1'b0;
  always @(*) begin
    LsuPlugin_logic_bus_cmd_ready = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_ready;
    if(when_Stream_l477_2) begin
      LsuPlugin_logic_bus_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l477_2 = (! LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid);
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid = LsuPlugin_logic_bus_cmd_rValid;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_write = LsuPlugin_logic_bus_cmd_rData_write;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_address = LsuPlugin_logic_bus_cmd_rData_address;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_data = LsuPlugin_logic_bus_cmd_rData_data;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_size = LsuPlugin_logic_bus_cmd_rData_size;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_mask = LsuPlugin_logic_bus_cmd_rData_mask;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_io = LsuPlugin_logic_bus_cmd_rData_io;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_fromHart = LsuPlugin_logic_bus_cmd_rData_fromHart;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_uopId = LsuPlugin_logic_bus_cmd_rData_uopId;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_ADR = (LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_address >>> 2'd3);
  assign LsuCachelessWishbonePlugin_logic_bridge_down_CTI = 3'b000;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_BTE = 2'b00;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_SEL = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_mask;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_WE = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_write;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_DAT_MOSI = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_payload_data;
  assign LsuCachelessWishbonePlugin_logic_bridge_cmdStage_ready = (LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid && (LsuCachelessWishbonePlugin_logic_bridge_down_ACK || LsuCachelessWishbonePlugin_logic_bridge_down_ERR));
  assign LsuCachelessWishbonePlugin_logic_bridge_down_CYC = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid;
  assign LsuCachelessWishbonePlugin_logic_bridge_down_STB = LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid;
  assign LsuPlugin_logic_bus_rsp_valid = (LsuCachelessWishbonePlugin_logic_bridge_cmdStage_valid && (LsuCachelessWishbonePlugin_logic_bridge_down_ACK || LsuCachelessWishbonePlugin_logic_bridge_down_ERR));
  assign LsuPlugin_logic_bus_rsp_payload_data = LsuCachelessWishbonePlugin_logic_bridge_down_DAT_MISO;
  assign LsuPlugin_logic_bus_rsp_payload_error = LsuCachelessWishbonePlugin_logic_bridge_down_ERR;
  assign LsuPlugin_logic_commitProbe_takeWhen_valid = (LsuPlugin_logic_commitProbe_valid && (! LsuPlugin_logic_commitProbe_payload_io));
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_pc = LsuPlugin_logic_commitProbe_payload_pc;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_address = LsuPlugin_logic_commitProbe_payload_address;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_load = LsuPlugin_logic_commitProbe_payload_load;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_store = LsuPlugin_logic_commitProbe_payload_store;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_trap = LsuPlugin_logic_commitProbe_payload_trap;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_io = LsuPlugin_logic_commitProbe_payload_io;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_prefetchFailed = LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  assign LsuPlugin_logic_commitProbe_takeWhen_payload_miss = LsuPlugin_logic_commitProbe_payload_miss;
  assign PrefetcherRptPlugin_logic_pip_node_0_valid = LsuPlugin_logic_commitProbe_takeWhen_valid;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_pc = LsuPlugin_logic_commitProbe_payload_pc;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_address = LsuPlugin_logic_commitProbe_payload_address;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_load = LsuPlugin_logic_commitProbe_payload_load;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_store = LsuPlugin_logic_commitProbe_payload_store;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_trap = LsuPlugin_logic_commitProbe_payload_trap;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_io = LsuPlugin_logic_commitProbe_payload_io;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_prefetchFailed = LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  assign PrefetcherRptPlugin_logic_pip_node_0_PROBE_miss = LsuPlugin_logic_commitProbe_payload_miss;
  assign PrefetcherRptPlugin_logic_storage_read_cmd_valid = PrefetcherRptPlugin_logic_pip_node_0_isFiring;
  assign PrefetcherRptPlugin_logic_storage_read_cmd_payload = PrefetcherRptPlugin_logic_pip_node_0_PROBE_pc[7 : 1];
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_valid = PrefetcherRptPlugin_logic_storage_write_valid;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_address = PrefetcherRptPlugin_logic_storage_write_payload_address;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_tag = PrefetcherRptPlugin_logic_storage_write_payload_data_tag;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_address = PrefetcherRptPlugin_logic_storage_write_payload_data_address;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_stride = PrefetcherRptPlugin_logic_storage_write_payload_data_stride;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_score = PrefetcherRptPlugin_logic_storage_write_payload_data_score;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_advance = PrefetcherRptPlugin_logic_storage_write_payload_data_advance;
  assign PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_missed = PrefetcherRptPlugin_logic_storage_write_payload_data_missed;
  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_tag = PrefetcherRptPlugin_logic_storage_read_rsp_tag;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_tag = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_tag;
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address = PrefetcherRptPlugin_logic_storage_read_rsp_address;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_address;
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_stride = PrefetcherRptPlugin_logic_storage_read_rsp_stride;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_stride = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_stride;
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_score = PrefetcherRptPlugin_logic_storage_read_rsp_score;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_score = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_score;
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_advance = PrefetcherRptPlugin_logic_storage_read_rsp_advance;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_advance = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_advance;
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_pip_node_1_ENTRY_missed = PrefetcherRptPlugin_logic_storage_read_rsp_missed;
    if(when_Prefetcher_l155) begin
      PrefetcherRptPlugin_logic_pip_node_1_ENTRY_missed = PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_missed;
    end
  end

  assign when_Prefetcher_l155 = (PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_valid && (PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_address == PrefetcherRptPlugin_logic_pip_node_1_PROBE_pc[7 : 1]));
  assign PrefetcherRptPlugin_logic_pip_node_1_TAG_HIT = (PrefetcherRptPlugin_logic_pip_node_1_ENTRY_tag == PrefetcherRptPlugin_logic_pip_node_1_PROBE_pc[22 : 8]);
  assign PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED = _zz_PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED[15:0];
  assign PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK = (_zz_PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK != 10'h0);
  assign _zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT = _zz__zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT;
  assign PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT = (($signed(_zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT_1) == $signed(PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride)) && (&{(_zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT[3] == PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride[11]),{(_zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT[2] == PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride[11]),{(_zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT[1] == PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride[11]),(_zz_PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT[0] == PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride[11])}}}));
  assign PrefetcherRptPlugin_logic_pip_node_2_STRIDE = PrefetcherRptPlugin_logic_pip_node_2_STRIDE_EXTENDED[11:0];
  always @(*) begin
    PrefetcherRptPlugin_logic_order_valid = PrefetcherRptPlugin_logic_onCtrl_unfiltred_valid;
    if(PrefetcherRptPlugin_logic_csr_disable) begin
      PrefetcherRptPlugin_logic_order_valid = 1'b0;
    end
  end

  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_ready = PrefetcherRptPlugin_logic_order_ready;
  assign PrefetcherRptPlugin_logic_order_payload_address = PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_address;
  assign PrefetcherRptPlugin_logic_order_payload_unique = PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_unique;
  assign PrefetcherRptPlugin_logic_order_payload_from = PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_from;
  assign PrefetcherRptPlugin_logic_order_payload_to = PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to;
  assign PrefetcherRptPlugin_logic_order_payload_stride = PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride;
  always @(*) begin
    PrefetcherRptPlugin_logic_onCtrl_add = 5'h0;
    if(!when_Prefetcher_l196) begin
      if(!when_Prefetcher_l208) begin
        if(PrefetcherRptPlugin_logic_pip_node_2_NEW_BLOCK) begin
          PrefetcherRptPlugin_logic_onCtrl_add = 5'h01;
        end
      end
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_onCtrl_sub = 5'h0;
    if(when_Prefetcher_l196) begin
      if(when_Prefetcher_l197) begin
        if(when_Prefetcher_l198) begin
          PrefetcherRptPlugin_logic_onCtrl_sub = 5'h02;
        end
      end
    end else begin
      if(when_Prefetcher_l208) begin
        PrefetcherRptPlugin_logic_onCtrl_sub = (PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score >>> 1);
      end
    end
  end

  assign _zz_when_UInt_l128 = ({1'b0,PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score} - {1'b0,PrefetcherRptPlugin_logic_onCtrl_sub});
  assign when_UInt_l128 = _zz_when_UInt_l128[5];
  always @(*) begin
    if(when_UInt_l128) begin
      _zz_PrefetcherRptPlugin_logic_onCtrl_score = 5'h0;
    end else begin
      _zz_PrefetcherRptPlugin_logic_onCtrl_score = _zz_when_UInt_l128[4 : 0];
    end
  end

  assign _zz_PrefetcherRptPlugin_logic_onCtrl_score_1 = ({1'b0,_zz_PrefetcherRptPlugin_logic_onCtrl_score} + {1'b0,PrefetcherRptPlugin_logic_onCtrl_add});
  assign when_UInt_l119_2 = (|_zz_PrefetcherRptPlugin_logic_onCtrl_score_1[5 : 5]);
  always @(*) begin
    if(when_UInt_l119_2) begin
      PrefetcherRptPlugin_logic_onCtrl_score = 5'h1f;
    end else begin
      PrefetcherRptPlugin_logic_onCtrl_score = _zz_PrefetcherRptPlugin_logic_onCtrl_score_1[4 : 0];
    end
  end

  assign _zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed = ({1'b0,((! PrefetcherRptPlugin_logic_pip_node_2_PROBE_miss) ? PrefetcherRptPlugin_logic_pip_node_2_ENTRY_advance : 3'b000)} - _zz__zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed);
  assign when_UInt_l128_1 = _zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed[3];
  always @(*) begin
    if(when_UInt_l128_1) begin
      PrefetcherRptPlugin_logic_onCtrl_advanceSubed = 3'b000;
    end else begin
      PrefetcherRptPlugin_logic_onCtrl_advanceSubed = _zz_PrefetcherRptPlugin_logic_onCtrl_advanceSubed[2 : 0];
    end
    if(!when_Prefetcher_l196) begin
      if(when_Prefetcher_l208) begin
        PrefetcherRptPlugin_logic_onCtrl_advanceSubed = 3'b000;
      end
    end
  end

  assign _zz_when_UInt_l128_1 = ({1'b0,PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score} - _zz__zz_when_UInt_l128_1);
  assign when_UInt_l128_2 = _zz_when_UInt_l128_1[5];
  always @(*) begin
    if(when_UInt_l128_2) begin
      _zz_PrefetcherRptPlugin_logic_onCtrl_advanceAllowed = 5'h0;
    end else begin
      _zz_PrefetcherRptPlugin_logic_onCtrl_advanceAllowed = _zz_when_UInt_l128_1[4 : 0];
    end
  end

  assign PrefetcherRptPlugin_logic_onCtrl_advanceAllowed = _zz_PrefetcherRptPlugin_logic_onCtrl_advanceAllowed;
  always @(*) begin
    PrefetcherRptPlugin_logic_onCtrl_orderAsk = 1'b0;
    if(!when_Prefetcher_l196) begin
      if(when_Prefetcher_l216) begin
        PrefetcherRptPlugin_logic_onCtrl_orderAsk = 1'b1;
      end
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_storage_write_valid = (PrefetcherRptPlugin_logic_pip_node_2_isFiring && (! PrefetcherRptPlugin_logic_pip_node_2_PROBE_prefetchFailed));
    if(PrefetcherRptPlugin_logic_csr_disable) begin
      PrefetcherRptPlugin_logic_storage_write_valid = 1'b0;
    end
  end

  assign PrefetcherRptPlugin_logic_storage_write_payload_address = PrefetcherRptPlugin_logic_pip_node_2_PROBE_pc[7 : 1];
  always @(*) begin
    PrefetcherRptPlugin_logic_storage_write_payload_data_tag = PrefetcherRptPlugin_logic_pip_node_2_ENTRY_tag;
    if(when_Prefetcher_l196) begin
      if(when_Prefetcher_l197) begin
        if(!when_Prefetcher_l198) begin
          PrefetcherRptPlugin_logic_storage_write_payload_data_tag = PrefetcherRptPlugin_logic_pip_node_2_PROBE_pc[22 : 8];
        end
      end
    end
  end

  assign PrefetcherRptPlugin_logic_storage_write_payload_data_address = (PrefetcherRptPlugin_logic_pip_node_2_PROBE_trap ? PrefetcherRptPlugin_logic_pip_node_2_ENTRY_address : _zz_PrefetcherRptPlugin_logic_storage_write_payload_data_address);
  always @(*) begin
    PrefetcherRptPlugin_logic_storage_write_payload_data_stride = ((PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score < 5'h03) ? PrefetcherRptPlugin_logic_pip_node_2_STRIDE : PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride);
    if(when_Prefetcher_l196) begin
      if(when_Prefetcher_l197) begin
        if(!when_Prefetcher_l198) begin
          PrefetcherRptPlugin_logic_storage_write_payload_data_stride = 12'h0;
        end
      end
    end
  end

  always @(*) begin
    PrefetcherRptPlugin_logic_storage_write_payload_data_score = PrefetcherRptPlugin_logic_onCtrl_score;
    if(when_Prefetcher_l196) begin
      if(when_Prefetcher_l197) begin
        if(!when_Prefetcher_l198) begin
          PrefetcherRptPlugin_logic_storage_write_payload_data_score = 5'h0;
        end
      end
    end
  end

  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_fire = (PrefetcherRptPlugin_logic_onCtrl_unfiltred_valid && PrefetcherRptPlugin_logic_onCtrl_unfiltred_ready);
  always @(*) begin
    PrefetcherRptPlugin_logic_storage_write_payload_data_advance = (PrefetcherRptPlugin_logic_onCtrl_unfiltred_fire ? PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to : PrefetcherRptPlugin_logic_onCtrl_advanceSubed);
    if(when_Prefetcher_l196) begin
      if(when_Prefetcher_l197) begin
        if(!when_Prefetcher_l198) begin
          PrefetcherRptPlugin_logic_storage_write_payload_data_advance = 3'b000;
        end
      end
    end
  end

  assign PrefetcherRptPlugin_logic_storage_write_payload_data_missed = (PrefetcherRptPlugin_logic_pip_node_2_PROBE_miss || (PrefetcherRptPlugin_logic_pip_node_2_ENTRY_missed && PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT));
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_valid = (((PrefetcherRptPlugin_logic_pip_node_2_isFiring && PrefetcherRptPlugin_logic_onCtrl_orderAsk) && (! PrefetcherRptPlugin_logic_pip_node_2_PROBE_prefetchFailed)) && PrefetcherRptPlugin_logic_storage_write_payload_data_missed);
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_address = PrefetcherRptPlugin_logic_pip_node_2_PROBE_address;
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_unique = PrefetcherRptPlugin_logic_pip_node_2_PROBE_store;
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_from = (PrefetcherRptPlugin_logic_onCtrl_advanceSubed + 3'b001);
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to = 3'b100;
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to = _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_to_1[2:0];
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride = 7'h40;
  assign _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_1 = 8'h40;
  assign PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride = (PrefetcherRptPlugin_logic_pip_node_2_STRIDE[11] ? _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_2 : _zz_PrefetcherRptPlugin_logic_onCtrl_unfiltred_payload_stride_5);
  assign when_Prefetcher_l196 = (! PrefetcherRptPlugin_logic_pip_node_2_TAG_HIT);
  assign when_Prefetcher_l197 = ($signed(PrefetcherRptPlugin_logic_pip_node_2_STRIDE) != $signed(12'h0));
  assign when_Prefetcher_l198 = (PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score != 5'h0);
  assign when_Prefetcher_l208 = (! PrefetcherRptPlugin_logic_pip_node_2_STRIDE_HIT);
  assign when_Prefetcher_l216 = ((PrefetcherRptPlugin_logic_onCtrl_advanceSubed < 3'b100) && (_zz_when_Prefetcher_l216 < PrefetcherRptPlugin_logic_onCtrl_advanceAllowed));
  assign PrefetcherRptPlugin_logic_pip_node_0_isFiring = (PrefetcherRptPlugin_logic_pip_node_0_isValid && PrefetcherRptPlugin_logic_pip_node_0_isReady);
  assign PrefetcherRptPlugin_logic_pip_node_0_isValid = PrefetcherRptPlugin_logic_pip_node_0_valid;
  assign PrefetcherRptPlugin_logic_pip_node_0_isReady = 1'b1;
  assign PrefetcherRptPlugin_logic_pip_node_1_isValid = PrefetcherRptPlugin_logic_pip_node_1_valid;
  assign PrefetcherRptPlugin_logic_pip_node_2_isFiring = (PrefetcherRptPlugin_logic_pip_node_2_isValid && PrefetcherRptPlugin_logic_pip_node_2_isReady);
  assign PrefetcherRptPlugin_logic_pip_node_2_isValid = PrefetcherRptPlugin_logic_pip_node_2_valid;
  assign PrefetcherRptPlugin_logic_pip_node_2_isReady = 1'b1;
  assign LsuPlugin_pmaBuilder_l1_addressBits = LsuPlugin_logic_onPma_cached_cmd_address;
  assign LsuPlugin_pmaBuilder_l1_argsBits = LsuPlugin_logic_onPma_cached_cmd_op;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io = ((LsuPlugin_pmaBuilder_l1_addressBits & 32'h0) == 32'h0);
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_l1_argsBits & 1'b0) == 1'b0));
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_hit = (LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit);
  assign LsuPlugin_logic_onPma_cached_rsp_fault = (! ((|((LsuPlugin_pmaBuilder_l1_addressBits & 32'h80000000) == 32'h80000000)) && (|LsuPlugin_pmaBuilder_l1_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_cached_rsp_io = (! _zz_LsuPlugin_logic_onPma_cached_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_io_addressBits = LsuPlugin_logic_onPma_io_cmd_address;
  assign LsuPlugin_pmaBuilder_io_argsBits = {LsuPlugin_logic_onPma_io_cmd_size,LsuPlugin_logic_onPma_io_cmd_op};
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_io_argsBits & 3'b000) == 3'b000));
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_hit = (LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault = ((LsuPlugin_pmaBuilder_io_addressBits & 32'h80000000) == 32'h80000000);
  assign LsuPlugin_logic_onPma_io_rsp_fault = (! ((|{_zz_LsuPlugin_logic_onPma_io_rsp_fault,((LsuPlugin_pmaBuilder_io_addressBits & 32'hf0000000) == 32'h10000000)}) && (|LsuPlugin_pmaBuilder_io_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_io_rsp_io = (! _zz_LsuPlugin_logic_onPma_io_rsp_io[0]);
  assign execute_ctrl2_COMPLETED_lane1_bypass = (execute_ctrl2_up_COMPLETED_lane1 || execute_ctrl2_down_COMPLETION_AT_2_lane1);
  assign execute_ctrl4_COMPLETED_lane1_bypass = (execute_ctrl4_up_COMPLETED_lane1 || execute_ctrl4_down_COMPLETION_AT_4_lane1);
  assign execute_lane1_api_hartsInflight[0] = (|{(execute_ctrl4_up_LANE_SEL_lane1 && 1'b1),{(execute_ctrl3_up_LANE_SEL_lane1 && 1'b1),{(execute_ctrl2_up_LANE_SEL_lane1 && 1'b1),(execute_ctrl1_up_LANE_SEL_lane1 && 1'b1)}}});
  assign _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX = FpuCmpPlugin_logic_ffwb_ats[0];
  assign execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX = (FpuCmpPlugin_logic_ffwb_flags_NX && _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX);
  assign execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF = (FpuCmpPlugin_logic_ffwb_flags_UF && _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX);
  assign execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF = (FpuCmpPlugin_logic_ffwb_flags_OF && _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX);
  assign execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ = (FpuCmpPlugin_logic_ffwb_flags_DZ && _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX);
  assign execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV = (FpuCmpPlugin_logic_ffwb_flags_NV && _zz_execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX);
  assign _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX = FpuF2iPlugin_logic_ffwb_ats[0];
  assign _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1 = FpuPackerPlugin_logic_flagsWb_ats[0];
  assign execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX = (execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX || ((FpuF2iPlugin_logic_ffwb_flags_NX && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX) || (FpuPackerPlugin_logic_flagsWb_flags_NX && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1)));
  assign execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_UF = (execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF || ((FpuF2iPlugin_logic_ffwb_flags_UF && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX) || (FpuPackerPlugin_logic_flagsWb_flags_UF && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1)));
  assign execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_OF = (execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF || ((FpuF2iPlugin_logic_ffwb_flags_OF && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX) || (FpuPackerPlugin_logic_flagsWb_flags_OF && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1)));
  assign execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_DZ = (execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ || ((FpuF2iPlugin_logic_ffwb_flags_DZ && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX) || (FpuPackerPlugin_logic_flagsWb_flags_DZ && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1)));
  assign execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NV = (execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV || ((FpuF2iPlugin_logic_ffwb_flags_NV && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX) || (FpuPackerPlugin_logic_flagsWb_flags_NV && _zz_execute_ctrl4_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_bypass_NX_1)));
  assign _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX = (execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_COMMIT_lane0);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX = (execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_0_UF = (execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_0_OF = (execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_0_DZ = (execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NV = (execute_ctrl4_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX);
  assign _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX = (|{((execute_ctrl11_up_LANE_SEL_lane0 && execute_ctrl11_up_COMMIT_lane0) && FpuPackerPlugin_logic_flagsWb_ats[4]),{((execute_ctrl8_up_LANE_SEL_lane0 && execute_ctrl8_up_COMMIT_lane0) && FpuPackerPlugin_logic_flagsWb_ats[3]),{((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_COMMIT_lane0) && FpuPackerPlugin_logic_flagsWb_ats[2]),((execute_ctrl7_up_LANE_SEL_lane0 && execute_ctrl7_up_COMMIT_lane0) && FpuPackerPlugin_logic_flagsWb_ats[1])}}});
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX = (FpuPackerPlugin_logic_flagsWb_flags_NX && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_1_UF = (FpuPackerPlugin_logic_flagsWb_flags_UF && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_1_OF = (FpuPackerPlugin_logic_flagsWb_flags_OF && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_1_DZ = (FpuPackerPlugin_logic_flagsWb_flags_DZ && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NV = (FpuPackerPlugin_logic_flagsWb_flags_NV && _zz_FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_flagsOr_NX = (FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NX || FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NX);
  assign FpuFlagsWritebackPlugin_logic_flagsOr_UF = (FpuFlagsWritebackPlugin_logic_afterCommit_0_0_UF || FpuFlagsWritebackPlugin_logic_afterCommit_0_1_UF);
  assign FpuFlagsWritebackPlugin_logic_flagsOr_OF = (FpuFlagsWritebackPlugin_logic_afterCommit_0_0_OF || FpuFlagsWritebackPlugin_logic_afterCommit_0_1_OF);
  assign FpuFlagsWritebackPlugin_logic_flagsOr_DZ = (FpuFlagsWritebackPlugin_logic_afterCommit_0_0_DZ || FpuFlagsWritebackPlugin_logic_afterCommit_0_1_DZ);
  assign FpuFlagsWritebackPlugin_logic_flagsOr_NV = (FpuFlagsWritebackPlugin_logic_afterCommit_0_0_NV || FpuFlagsWritebackPlugin_logic_afterCommit_0_1_NV);
  assign execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0) == $signed(execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0));
  assign execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0 != execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign late0_BranchPlugin_logic_alu_expectedMsb = 1'b0;
  assign execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l245_3 = execute_ctrl4_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l245_3)
      3'b000 : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl4_down_late0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 ? execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0 != execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_needFix = ((late0_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 && execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_late0_BranchPlugin_SEL_lane0) && late0_BranchPlugin_logic_jumpLogic_needFix);
  assign late0_BranchPlugin_logic_jumpLogic_history_slice = execute_ctrl4_down_PC_lane0[2 : 1];
  assign late0_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l213_6 = ((late0_BranchPlugin_logic_jumpLogic_history_slice < 2'b00) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[0]);
  assign when_BranchPlugin_l213_7 = ((late0_BranchPlugin_logic_jumpLogic_history_slice < 2'b01) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[1]);
  assign when_BranchPlugin_l213_8 = ((late0_BranchPlugin_logic_jumpLogic_history_slice < 2'b10) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[2]);
  assign when_BranchPlugin_l218_2 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign late0_BranchPlugin_logic_jumpLogic_history_next = late0_BranchPlugin_logic_jumpLogic_history_shifter_4;
  assign late0_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  assign late0_BranchPlugin_logic_pcPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign late0_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign late0_BranchPlugin_logic_pcPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_historyPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_historyPort_payload_history = late0_BranchPlugin_logic_jumpLogic_history_next;
  assign late0_BranchPlugin_logic_historyPort_payload_age = execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_flushPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign late0_BranchPlugin_logic_flushPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0 : 0] != 1'b0) && execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign late0_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == 5'h05),(execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign late0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl4_down_Decode_UOP_lane0[19 : 15] == 5'h05),(execute_ctrl4_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign late0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == execute_ctrl4_down_Decode_UOP_lane0[19 : 15]);
  assign late0_BranchPlugin_logic_jumpLogic_learn_valid = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && (|{execute_ctrl4_down_late0_BranchPlugin_SEL_lane0,execute_ctrl4_down_early0_BranchPlugin_SEL_lane0}));
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_taken = execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 || execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0) && late0_BranchPlugin_logic_jumpLogic_rdLink);
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 && (((! late0_BranchPlugin_logic_jumpLogic_rdLink) && late0_BranchPlugin_logic_jumpLogic_rs1Link) || ((late0_BranchPlugin_logic_jumpLogic_rdLink && late0_BranchPlugin_logic_jumpLogic_rs1Link) && (! late0_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_needFix;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_history = late0_BranchPlugin_logic_jumpLogic_history_fetched;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign late0_BranchPlugin_logic_wb_valid = execute_ctrl4_down_late0_BranchPlugin_SEL_lane0;
  assign late0_BranchPlugin_logic_wb_payload = execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1 = ($signed(execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1) == $signed(execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1));
  assign execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 = (execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1 != execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1);
  assign late1_BranchPlugin_logic_alu_expectedMsb = 1'b0;
  assign execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1 = ((execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l245_4 = execute_ctrl4_down_Decode_UOP_lane1[14 : 12];
  always @(*) begin
    casez(switch_Misc_l245_4)
      3'b000 : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1;
      end
      3'b001 : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1);
      end
      3'b1?1 : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! execute_ctrl4_down_late1_SrcPlugin_LESS_lane1);
      end
      default : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
      end
    endcase
  end

  assign execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = _zz_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  assign execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1 = (execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 ? execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 : execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1 != execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_needFix = ((late1_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 && execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1)) || execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_down_late1_BranchPlugin_SEL_lane1) && late1_BranchPlugin_logic_jumpLogic_needFix);
  assign late1_BranchPlugin_logic_jumpLogic_history_slice = execute_ctrl4_down_PC_lane1[2 : 1];
  assign late1_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  assign when_BranchPlugin_l213_9 = ((late1_BranchPlugin_logic_jumpLogic_history_slice < 2'b00) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[0]);
  assign when_BranchPlugin_l213_10 = ((late1_BranchPlugin_logic_jumpLogic_history_slice < 2'b01) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[1]);
  assign when_BranchPlugin_l213_11 = ((late1_BranchPlugin_logic_jumpLogic_history_slice < 2'b10) && execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[2]);
  assign when_BranchPlugin_l218_3 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign late1_BranchPlugin_logic_jumpLogic_history_next = late1_BranchPlugin_logic_jumpLogic_history_shifter_4;
  assign late1_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  assign late1_BranchPlugin_logic_pcPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  assign late1_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  assign late1_BranchPlugin_logic_pcPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_historyPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_historyPort_payload_history = late1_BranchPlugin_logic_jumpLogic_history_next;
  assign late1_BranchPlugin_logic_historyPort_payload_age = execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_flushPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign late1_BranchPlugin_logic_flushPort_payload_laneAge = execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1 = ((execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0 : 0] != 1'b0) && execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR);
  assign late1_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == 5'h05),(execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == 5'h01)});
  assign late1_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl4_down_Decode_UOP_lane1[19 : 15] == 5'h05),(execute_ctrl4_down_Decode_UOP_lane1[19 : 15] == 5'h01)});
  assign late1_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == execute_ctrl4_down_Decode_UOP_lane1[19 : 15]);
  assign late1_BranchPlugin_logic_jumpLogic_learn_valid = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_upIsCancel)) && (|{execute_ctrl4_down_late1_BranchPlugin_SEL_lane1,execute_ctrl4_down_early1_BranchPlugin_SEL_lane1}));
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_taken = execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 || execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1) && late1_BranchPlugin_logic_jumpLogic_rdLink);
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 && (((! late1_BranchPlugin_logic_jumpLogic_rdLink) && late1_BranchPlugin_logic_jumpLogic_rs1Link) || ((late1_BranchPlugin_logic_jumpLogic_rdLink && late1_BranchPlugin_logic_jumpLogic_rs1Link) && (! late1_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_needFix;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_history = late1_BranchPlugin_logic_jumpLogic_history_fetched;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign late1_BranchPlugin_logic_wb_valid = execute_ctrl4_down_late1_BranchPlugin_SEL_lane1;
  assign late1_BranchPlugin_logic_wb_payload = execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign execute_ctrl4_COMPLETED_lane0_bypass = (execute_ctrl4_up_COMPLETED_lane0 || execute_ctrl4_down_COMPLETION_AT_4_lane0);
  assign execute_ctrl7_COMPLETED_lane0_bypass = (execute_ctrl7_up_COMPLETED_lane0 || execute_ctrl7_down_COMPLETION_AT_7_lane0);
  assign execute_ctrl11_COMPLETED_lane0_bypass = (execute_ctrl11_up_COMPLETED_lane0 || execute_ctrl11_down_COMPLETION_AT_11_lane0);
  assign execute_ctrl3_COMPLETED_lane0_bypass = (execute_ctrl3_up_COMPLETED_lane0 || execute_ctrl3_down_COMPLETION_AT_3_lane0);
  assign execute_ctrl5_COMPLETED_lane0_bypass = (execute_ctrl5_up_COMPLETED_lane0 || execute_ctrl5_down_COMPLETION_AT_5_lane0);
  assign execute_ctrl8_COMPLETED_lane0_bypass = (execute_ctrl8_up_COMPLETED_lane0 || execute_ctrl8_down_COMPLETION_AT_8_lane0);
  assign execute_ctrl2_COMPLETED_lane0_bypass = (execute_ctrl2_up_COMPLETED_lane0 || execute_ctrl2_down_COMPLETION_AT_2_lane0);
  assign execute_lane0_api_hartsInflight[0] = (|{((execute_ctrl11_up_LANE_SEL_lane0 && (! execute_ctrl11_down_COMPLETED_lane0)) && 1'b1),{((execute_ctrl10_up_LANE_SEL_lane0 && (! execute_ctrl10_down_COMPLETED_lane0)) && 1'b1),{((execute_ctrl9_up_LANE_SEL_lane0 && _zz_execute_lane0_api_hartsInflight) && 1'b1),{(_zz_execute_lane0_api_hartsInflight_1 && _zz_execute_lane0_api_hartsInflight_2),{_zz_execute_lane0_api_hartsInflight_3,{_zz_execute_lane0_api_hartsInflight_4,_zz_execute_lane0_api_hartsInflight_5}}}}}});
  assign _zz_CsrRamPlugin_csrMapper_ramAddress = CsrAccessPlugin_bus_decode_address;
  assign CsrRamPlugin_csrMapper_ramAddress = {(|{((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h002) == 12'h002),((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h040) == 12'h0)}),(|((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h003) == 12'h001))};
  always @(*) begin
    CsrRamPlugin_csrMapper_withRead = 1'b0;
    if(when_CsrAccessPlugin_l252) begin
      CsrRamPlugin_csrMapper_withRead = 1'b1;
    end
  end

  assign CsrRamPlugin_csrMapper_read_valid = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_api_holdRead));
  assign CsrRamPlugin_csrMapper_read_address = CsrRamPlugin_csrMapper_ramAddress;
  assign when_CsrRamPlugin_l85 = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_csrMapper_read_ready));
  always @(*) begin
    CsrRamPlugin_csrMapper_doWrite = 1'b0;
    if(when_CsrAccessPlugin_l343_2) begin
      CsrRamPlugin_csrMapper_doWrite = 1'b1;
    end
  end

  assign when_CsrRamPlugin_l92 = (CsrRamPlugin_csrMapper_write_valid && CsrRamPlugin_csrMapper_write_ready);
  assign CsrRamPlugin_csrMapper_write_valid = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_api_holdWrite));
  assign CsrRamPlugin_csrMapper_write_address = CsrRamPlugin_csrMapper_ramAddress;
  assign CsrRamPlugin_csrMapper_write_data = CsrAccessPlugin_bus_write_bits;
  assign when_CsrRamPlugin_l96 = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_csrMapper_write_ready));
  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_learn_ready = LearnPlugin_logic_buffered_0_ready;
    if(when_Stream_l477_3) begin
      late0_BranchPlugin_logic_jumpLogic_learn_ready = 1'b1;
    end
  end

  assign when_Stream_l477_3 = (! LearnPlugin_logic_buffered_0_valid);
  assign LearnPlugin_logic_buffered_0_valid = late0_BranchPlugin_logic_jumpLogic_learn_rValid;
  assign LearnPlugin_logic_buffered_0_payload_pcOnLastSlice = late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  assign LearnPlugin_logic_buffered_0_payload_pcTarget = late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  assign LearnPlugin_logic_buffered_0_payload_taken = late0_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  assign LearnPlugin_logic_buffered_0_payload_isBranch = late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  assign LearnPlugin_logic_buffered_0_payload_isPush = late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  assign LearnPlugin_logic_buffered_0_payload_isPop = late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  assign LearnPlugin_logic_buffered_0_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  assign LearnPlugin_logic_buffered_0_payload_badPredictedTarget = late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  assign LearnPlugin_logic_buffered_0_payload_history = late0_BranchPlugin_logic_jumpLogic_learn_rData_history;
  assign LearnPlugin_logic_buffered_0_payload_uopId = late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_learn_ready = LearnPlugin_logic_buffered_1_ready;
    if(when_Stream_l477_4) begin
      late1_BranchPlugin_logic_jumpLogic_learn_ready = 1'b1;
    end
  end

  assign when_Stream_l477_4 = (! LearnPlugin_logic_buffered_1_valid);
  assign LearnPlugin_logic_buffered_1_valid = late1_BranchPlugin_logic_jumpLogic_learn_rValid;
  assign LearnPlugin_logic_buffered_1_payload_pcOnLastSlice = late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  assign LearnPlugin_logic_buffered_1_payload_pcTarget = late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  assign LearnPlugin_logic_buffered_1_payload_taken = late1_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  assign LearnPlugin_logic_buffered_1_payload_isBranch = late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  assign LearnPlugin_logic_buffered_1_payload_isPush = late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  assign LearnPlugin_logic_buffered_1_payload_isPop = late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  assign LearnPlugin_logic_buffered_1_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  assign LearnPlugin_logic_buffered_1_payload_badPredictedTarget = late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  assign LearnPlugin_logic_buffered_1_payload_history = late1_BranchPlugin_logic_jumpLogic_learn_rData_history;
  assign LearnPlugin_logic_buffered_1_payload_uopId = late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  assign LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_buffered_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign LearnPlugin_logic_buffered_0_ready = streamArbiter_5_io_inputs_0_ready;
  assign LearnPlugin_logic_buffered_1_ready = streamArbiter_5_io_inputs_1_ready;
  assign LearnPlugin_logic_arbitrated_valid = streamArbiter_5_io_output_valid;
  assign LearnPlugin_logic_arbitrated_payload_pcOnLastSlice = streamArbiter_5_io_output_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_payload_pcTarget = streamArbiter_5_io_output_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_payload_taken = streamArbiter_5_io_output_payload_taken;
  assign LearnPlugin_logic_arbitrated_payload_isBranch = streamArbiter_5_io_output_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_payload_isPush = streamArbiter_5_io_output_payload_isPush;
  assign LearnPlugin_logic_arbitrated_payload_isPop = streamArbiter_5_io_output_payload_isPop;
  assign LearnPlugin_logic_arbitrated_payload_wasWrong = streamArbiter_5_io_output_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_payload_badPredictedTarget = streamArbiter_5_io_output_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_payload_history = streamArbiter_5_io_output_payload_history;
  assign LearnPlugin_logic_arbitrated_payload_uopId = streamArbiter_5_io_output_payload_uopId;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = streamArbiter_5_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign LearnPlugin_logic_arbitrated_ready = 1'b1;
  assign LearnPlugin_logic_arbitrated_toFlow_valid = LearnPlugin_logic_arbitrated_valid;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget = LearnPlugin_logic_arbitrated_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_taken = LearnPlugin_logic_arbitrated_payload_taken;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isBranch = LearnPlugin_logic_arbitrated_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPush = LearnPlugin_logic_arbitrated_payload_isPush;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPop = LearnPlugin_logic_arbitrated_payload_isPop;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong = LearnPlugin_logic_arbitrated_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_history = LearnPlugin_logic_arbitrated_payload_history;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_uopId = LearnPlugin_logic_arbitrated_payload_uopId;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign LearnPlugin_logic_learn_valid = LearnPlugin_logic_arbitrated_toFlow_valid;
  assign LearnPlugin_logic_learn_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  assign LearnPlugin_logic_learn_payload_pcTarget = LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  assign LearnPlugin_logic_learn_payload_taken = LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  assign LearnPlugin_logic_learn_payload_isBranch = LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  assign LearnPlugin_logic_learn_payload_isPush = LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  assign LearnPlugin_logic_learn_payload_isPop = LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  assign LearnPlugin_logic_learn_payload_wasWrong = LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  assign LearnPlugin_logic_learn_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  assign LearnPlugin_logic_learn_payload_history = LearnPlugin_logic_arbitrated_toFlow_payload_history;
  assign LearnPlugin_logic_learn_payload_uopId = LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign when_DecoderPlugin_l143 = (decode_ctrls_1_up_isMoving && 1'b1);
  assign DecoderPlugin_logic_interrupt_async = PrivilegedPlugin_logic_harts_0_int_pending;
  assign when_DecoderPlugin_l151 = (((! decode_ctrls_1_up_valid) || decode_ctrls_1_up_ready) || decode_ctrls_1_up_isCanceling);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000060) == 32'h00000040);
  assign decode_ctrls_1_down_RS1_ENABLE_0 = _zz_decode_ctrls_1_down_RS1_ENABLE_0[0];
  assign _zz_decode_ctrls_1_down_RD_RFID_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h80000060) == 32'h00000040);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000070) == 32'h00000040);
  assign decode_ctrls_1_down_RS1_RFID_0 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0,{_zz_decode_ctrls_1_down_RD_RFID_0,((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h10000060) == 32'h00000040)}});
  assign decode_ctrls_1_down_RS1_PHYS_0 = _zz_decode_ctrls_1_down_RS1_PHYS_0[4 : 0];
  assign decode_ctrls_1_down_RS2_ENABLE_0 = _zz_decode_ctrls_1_down_RS2_ENABLE_0[0];
  assign decode_ctrls_1_down_RS2_RFID_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000020) == 32'h0),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000000c) == 32'h00000004)});
  assign decode_ctrls_1_down_RS2_PHYS_0 = _zz_decode_ctrls_1_down_RS2_PHYS_0[4 : 0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000014) == 32'h00000014);
  always @(*) begin
    decode_ctrls_1_down_RD_ENABLE_0 = _zz_decode_ctrls_1_down_RD_ENABLE_0[0];
    if(when_DecoderPlugin_l247) begin
      decode_ctrls_1_down_RD_ENABLE_0 = 1'b0;
    end
  end

  assign decode_ctrls_1_down_RD_RFID_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h10000060) == 32'h10000040),{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0,{_zz_decode_ctrls_1_down_RD_RFID_0,((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000034) == 32'h00000004)}}});
  assign decode_ctrls_1_down_RD_PHYS_0 = _zz_decode_ctrls_1_down_RD_PHYS_0[4 : 0];
  assign decode_ctrls_1_down_RS3_ENABLE_0 = _zz_decode_ctrls_1_down_RS3_ENABLE_0[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0) == 32'h0);
  assign decode_ctrls_1_down_RS3_RFID_0 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign decode_ctrls_1_down_RS3_PHYS_0 = _zz_decode_ctrls_1_down_RS3_PHYS_0[4 : 0];
  always @(*) begin
    decode_ctrls_1_down_Decode_LEGAL_0 = ((|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005f) == 32'h00000017),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h04000073) == 32'h00000043),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0) == 32'h0000006f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_1 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_2),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_3,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_4,_zz_decode_ctrls_1_down_Decode_LEGAL_0_5}}}}}}) && (! decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0));
    if(DecoderPlugin_logic_laneLogic_0_fp_triggered) begin
      decode_ctrls_1_down_Decode_LEGAL_0 = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_fp_instRm = decode_ctrls_1_down_Decode_UOP_0[14 : 12];
  assign DecoderPlugin_logic_laneLogic_0_fp_rm = ((DecoderPlugin_logic_laneLogic_0_fp_instRm == 3'b111) ? FpuCsrPlugin_api_rm : DecoderPlugin_logic_laneLogic_0_fp_instRm);
  assign DecoderPlugin_logic_laneLogic_0_fp_triggered = ((decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 && (! PrivilegedPlugin_api_harts_0_fpuEnable)) || (decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 && (3'b101 <= DecoderPlugin_logic_laneLogic_0_fp_rm)));
  assign DecoderPlugin_logic_laneLogic_0_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l229) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_valid = ((! decode_ctrls_1_up_TRAP_0) || DecoderPlugin_logic_laneLogic_0_interruptPending);
      if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval = decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge = 2'b00;
  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg = 2'b00;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000070) == 32'h00000060);
  assign DecoderPlugin_logic_laneLogic_0_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_0_fixer_doIt = (decode_ctrls_1_up_LANE_SEL_0 && ((decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 && (! DecoderPlugin_logic_laneLogic_0_fixer_isJb)) || decode_ctrls_1_down_Prediction_ALIGN_REDO_0));
  assign when_CtrlLaneApi_l50_2 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_0_completionPort_valid = ((decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0) && (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext)));
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l229 = (decode_ctrls_1_up_LANE_SEL_0 && (((! decode_ctrls_1_down_Decode_LEGAL_0) || DecoderPlugin_logic_laneLogic_0_interruptPending) || DecoderPlugin_logic_laneLogic_0_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_0_flushPort_valid = (decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0);
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge = 1'b0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l247 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7] == 5'h0) && (|(decode_ctrls_1_down_RD_RFID_0 == 1'b0)));
  assign decode_ctrls_1_down_Decode_UOP_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0;
  assign DecoderPlugin_logic_laneLogic_0_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign decode_ctrls_1_down_Decode_UOP_ID_0 = (DecoderPlugin_logic_laneLogic_0_uopIdBase + 16'h0);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000060) == 32'h00000040);
  assign decode_ctrls_1_down_RS1_ENABLE_1 = _zz_decode_ctrls_1_down_RS1_ENABLE_1[0];
  assign _zz_decode_ctrls_1_down_RD_RFID_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h80000060) == 32'h00000040);
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000070) == 32'h00000040);
  assign decode_ctrls_1_down_RS1_RFID_1 = (|{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1,{_zz_decode_ctrls_1_down_RD_RFID_1,((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h10000060) == 32'h00000040)}});
  assign decode_ctrls_1_down_RS1_PHYS_1 = _zz_decode_ctrls_1_down_RS1_PHYS_1[4 : 0];
  assign decode_ctrls_1_down_RS2_ENABLE_1 = _zz_decode_ctrls_1_down_RS2_ENABLE_1[0];
  assign decode_ctrls_1_down_RS2_RFID_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000020) == 32'h0),((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000000c) == 32'h00000004)});
  assign decode_ctrls_1_down_RS2_PHYS_1 = _zz_decode_ctrls_1_down_RS2_PHYS_1[4 : 0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000014) == 32'h00000014);
  always @(*) begin
    decode_ctrls_1_down_RD_ENABLE_1 = _zz_decode_ctrls_1_down_RD_ENABLE_1[0];
    if(when_DecoderPlugin_l247_1) begin
      decode_ctrls_1_down_RD_ENABLE_1 = 1'b0;
    end
  end

  assign decode_ctrls_1_down_RD_RFID_1 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h10000060) == 32'h10000040),{_zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1,{_zz_decode_ctrls_1_down_RD_RFID_1,((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000034) == 32'h00000004)}}});
  assign decode_ctrls_1_down_RD_PHYS_1 = _zz_decode_ctrls_1_down_RD_PHYS_1[4 : 0];
  assign decode_ctrls_1_down_RS3_ENABLE_1 = _zz_decode_ctrls_1_down_RS3_ENABLE_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0) == 32'h0);
  assign decode_ctrls_1_down_RS3_RFID_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign decode_ctrls_1_down_RS3_PHYS_1 = _zz_decode_ctrls_1_down_RS3_PHYS_1[4 : 0];
  always @(*) begin
    decode_ctrls_1_down_Decode_LEGAL_1 = ((|{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000005f) == 32'h00000017),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h04000073) == 32'h00000043),{((decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_decode_ctrls_1_down_Decode_LEGAL_1) == 32'h0000006f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_1_1 == _zz_decode_ctrls_1_down_Decode_LEGAL_1_2),{_zz_decode_ctrls_1_down_Decode_LEGAL_1_3,{_zz_decode_ctrls_1_down_Decode_LEGAL_1_4,_zz_decode_ctrls_1_down_Decode_LEGAL_1_5}}}}}}) && (! decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1));
    if(DecoderPlugin_logic_laneLogic_1_fp_triggered) begin
      decode_ctrls_1_down_Decode_LEGAL_1 = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_1_fp_instRm = decode_ctrls_1_down_Decode_UOP_1[14 : 12];
  assign DecoderPlugin_logic_laneLogic_1_fp_rm = ((DecoderPlugin_logic_laneLogic_1_fp_instRm == 3'b111) ? FpuCsrPlugin_api_rm : DecoderPlugin_logic_laneLogic_1_fp_instRm);
  assign DecoderPlugin_logic_laneLogic_1_fp_triggered = ((decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1 && (! PrivilegedPlugin_api_harts_0_fpuEnable)) || (decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1 && (3'b101 <= DecoderPlugin_logic_laneLogic_1_fp_rm)));
  assign DecoderPlugin_logic_laneLogic_1_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l229_1) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_valid = ((! decode_ctrls_1_up_TRAP_1) || DecoderPlugin_logic_laneLogic_1_interruptPending);
      if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_1_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_1_interruptPending) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval = decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1;
  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_1_interruptPending) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge = 2'b01;
  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg = 2'b00;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000070) == 32'h00000060);
  assign DecoderPlugin_logic_laneLogic_1_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_1_fixer_doIt = (decode_ctrls_1_up_LANE_SEL_1 && ((decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1 && (! DecoderPlugin_logic_laneLogic_1_fixer_isJb)) || decode_ctrls_1_down_Prediction_ALIGN_REDO_1));
  assign when_CtrlLaneApi_l50_3 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane1_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_1_completionPort_valid = ((decode_ctrls_1_up_LANE_SEL_1 && decode_ctrls_1_down_TRAP_1) && (decode_ctrls_1_up_LANE_SEL_1 && (! decode_ctrls_1_up_LANE_SEL_1_regNext)));
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l229_1 = (decode_ctrls_1_up_LANE_SEL_1 && (((! decode_ctrls_1_down_Decode_LEGAL_1) || DecoderPlugin_logic_laneLogic_1_interruptPending) || DecoderPlugin_logic_laneLogic_1_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_1_flushPort_valid = (decode_ctrls_1_up_LANE_SEL_1 && decode_ctrls_1_down_TRAP_1);
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge = 1'b1;
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l247_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1[11 : 7] == 5'h0) && (|(decode_ctrls_1_down_RD_RFID_1 == 1'b0)));
  assign decode_ctrls_1_down_Decode_UOP_1 = decode_ctrls_1_down_Decode_INSTRUCTION_1;
  assign DecoderPlugin_logic_laneLogic_1_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign decode_ctrls_1_down_Decode_UOP_ID_1 = (DecoderPlugin_logic_laneLogic_1_uopIdBase + 16'h0001);
  assign DispatchPlugin_logic_trapPendings[0] = (|(DispatchPlugin_logic_slots_0_ctx_valid && DispatchPlugin_logic_slots_0_ctx_hm_TRAP));
  assign DispatchPlugin_logic_candidates_0_moving = (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_candidates_0_fire) || DispatchPlugin_logic_candidates_0_cancel);
  assign DispatchPlugin_logic_candidates_1_moving = (((! DispatchPlugin_logic_candidates_1_ctx_valid) || DispatchPlugin_logic_candidates_1_fire) || DispatchPlugin_logic_candidates_1_cancel);
  assign DispatchPlugin_logic_candidates_2_moving = (((! DispatchPlugin_logic_candidates_2_ctx_valid) || DispatchPlugin_logic_candidates_2_fire) || DispatchPlugin_logic_candidates_2_cancel);
  assign DispatchPlugin_logic_candidates_0_age = 1'b0;
  assign DispatchPlugin_logic_candidates_1_age = _zz_DispatchPlugin_logic_candidates_1_age;
  assign DispatchPlugin_logic_candidates_2_age = _zz_DispatchPlugin_logic_candidates_2_age[0:0];
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5),(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_6 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_7)}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_2_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE && 1'b0);
  always @(*) begin
    DispatchPlugin_logic_candidates_0_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_0_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_0_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_0_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard}});
  end

  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_9,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_12}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_9,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_12}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE && (|{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_1) && (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID)) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_3) && (! execute_ctrl8_down_BYPASSED_AT_9_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_9,_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_2_hazard_12}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_2_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_2_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_2_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE && 1'b0);
  always @(*) begin
    DispatchPlugin_logic_candidates_1_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_1_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_1_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_1_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard}});
  end

  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_9,_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_12}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_9,_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_12}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID)) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_1) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID)) && (! execute_ctrl8_down_BYPASSED_AT_9_lane0)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_3) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_7,_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_2_hazard_10}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_2_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_2_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_2_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && 1'b0);
  always @(*) begin
    DispatchPlugin_logic_candidates_2_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_2_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_2_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard}});
    DispatchPlugin_logic_candidates_2_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_2_hazard,{DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard}});
  end

  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_7,_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_10}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (execute_ctrl2_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1) && (execute_ctrl1_up_RD_RFID_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID)) && (! execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_7,_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_10}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (execute_ctrl9_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID)) && (! execute_ctrl9_down_BYPASSED_AT_10_lane0)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_1) && (execute_ctrl8_up_RD_RFID_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID)) && (! execute_ctrl8_down_BYPASSED_AT_9_lane0)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_3) && (! execute_ctrl7_down_BYPASSED_AT_8_lane0)),{(_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_5),{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_6,{_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_7,_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_2_hazard_10}}}}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_2_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_2_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && 1'b0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_0_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_0_onLl_1_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_0_onLl_2_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_0_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_0_checks_0_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_2_checks_0_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_0_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_1_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_0_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_1_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_2_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl7_up_LANE_SEL_lane0) && execute_ctrl7_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_3_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_0_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_1_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl2_up_LANE_SEL_lane0) && execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_2_hit = ((DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl6_up_LANE_SEL_lane0) && execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_hit = (|{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_2_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_1_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_6_checks_0_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_3_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_2_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_1_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_5_checks_0_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_1_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_3_checks_0_hit,{DispatchPlugin_logic_reservationChecker_0_onLl_1_res_2_checks_0_hit,DispatchPlugin_logic_reservationChecker_0_onLl_1_res_0_checks_0_hit}}}}}}}}}});
  assign DispatchPlugin_logic_reservationChecker_0_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_0_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_1_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_1_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_1_onLl_0_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_1_onLl_1_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_1_onLl_2_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_1_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_0_checks_0_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_2_checks_0_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_0_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_1_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_0_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_1_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_2_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl7_up_LANE_SEL_lane0) && execute_ctrl7_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_3_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_0_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_1_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl2_up_LANE_SEL_lane0) && execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_2_hit = ((DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl6_up_LANE_SEL_lane0) && execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_hit = (|{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_2_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_1_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_6_checks_0_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_3_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_2_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_1_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_5_checks_0_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_1_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_3_checks_0_hit,{DispatchPlugin_logic_reservationChecker_1_onLl_1_res_2_checks_0_hit,DispatchPlugin_logic_reservationChecker_1_onLl_1_res_0_checks_0_hit}}}}}}}}}});
  assign DispatchPlugin_logic_reservationChecker_1_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_1_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_2_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_2_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_2_onLl_0_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_2_onLl_1_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_2_onLl_2_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_2_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_0_checks_0_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_2_checks_0_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_0_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_1_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_0_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_1_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_2_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl7_up_LANE_SEL_lane0) && execute_ctrl7_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_3_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 && execute_ctrl1_up_LANE_SEL_lane0) && execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_0_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl3_up_LANE_SEL_lane0) && execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_1_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl2_up_LANE_SEL_lane0) && execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_2_hit = ((DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 && execute_ctrl6_up_LANE_SEL_lane0) && execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0);
  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_hit = (|{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_2_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_1_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_6_checks_0_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_3_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_2_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_1_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_5_checks_0_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_1_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_3_checks_0_hit,{DispatchPlugin_logic_reservationChecker_2_onLl_1_res_2_checks_0_hit,DispatchPlugin_logic_reservationChecker_2_onLl_1_res_0_checks_0_hit}}}}}}}}}});
  assign DispatchPlugin_logic_reservationChecker_2_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_2_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_0_oldersHazard = 1'b0;
  assign DispatchPlugin_logic_candidates_0_flushHazards = ((|{DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_0_oldersHazard));
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_1_oldersHazard = (|(DispatchPlugin_logic_candidates_0_ctx_valid && DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH));
  assign DispatchPlugin_logic_candidates_1_flushHazards = ((|{DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_1_oldersHazard));
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_2_oldersHazard = (|{(DispatchPlugin_logic_candidates_1_ctx_valid && DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH),(DispatchPlugin_logic_candidates_0_ctx_valid && DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH)});
  assign DispatchPlugin_logic_candidates_2_flushHazards = ((|{DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_2_oldersHazard));
  assign DispatchPlugin_logic_fenceChecker_olderInflights = (|{execute_lane1_api_hartsInflight[0],execute_lane0_api_hartsInflight[0]});
  assign DispatchPlugin_logic_candidates_0_fenceOlderHazards = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || 1'b0));
  assign DispatchPlugin_logic_candidates_1_fenceOlderHazards = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || (|(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1))));
  assign DispatchPlugin_logic_candidates_2_fenceOlderHazards = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || (|{(DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1),(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1)})));
  always @(*) begin
    decode_ctrls_1_down_ready = 1'b1;
    if(when_DispatchPlugin_l368) begin
      decode_ctrls_1_down_ready = 1'b0;
    end
    if(when_DispatchPlugin_l368_1) begin
      decode_ctrls_1_down_ready = 1'b0;
    end
    if(DispatchPlugin_logic_slotsFeeds_doIt) begin
      decode_ctrls_1_down_ready = 1'b1;
    end
  end

  assign DispatchPlugin_logic_feeds_0_sending = DispatchPlugin_logic_candidates_1_fire;
  assign DispatchPlugin_logic_candidates_1_cancel = decode_ctrls_1_lane0_upIsCancel;
  assign DispatchPlugin_logic_candidates_1_ctx_valid = ((decode_ctrls_1_up_isValid && decode_ctrls_1_up_LANE_SEL_0) && (! DispatchPlugin_logic_feeds_0_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_1_ctx_laneLayerHits = {decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0,{decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0,decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0}}};
    if(decode_ctrls_1_down_TRAP_0) begin
      DispatchPlugin_logic_candidates_1_ctx_laneLayerHits = 4'b0010;
    end
  end

  assign DispatchPlugin_logic_candidates_1_ctx_uop = decode_ctrls_1_down_Decode_UOP_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY = decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER = decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH = decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 = decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 = decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_PC = decode_ctrls_1_down_PC_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_TRAP = decode_ctrls_1_down_TRAP_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE = decode_ctrls_1_down_RS1_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID = decode_ctrls_1_down_RS1_RFID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS = decode_ctrls_1_down_RS1_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE = decode_ctrls_1_down_RS2_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID = decode_ctrls_1_down_RS2_RFID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS = decode_ctrls_1_down_RS2_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE = decode_ctrls_1_down_RD_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID = decode_ctrls_1_down_RD_RFID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS = decode_ctrls_1_down_RD_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE = decode_ctrls_1_down_RS3_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID = decode_ctrls_1_down_RS3_RFID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS = decode_ctrls_1_down_RS3_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  assign when_DispatchPlugin_l368 = ((decode_ctrls_1_up_LANE_SEL_0 && (! DispatchPlugin_logic_feeds_0_sent)) && (! DispatchPlugin_logic_candidates_1_fire));
  assign DispatchPlugin_logic_feeds_1_sending = DispatchPlugin_logic_candidates_2_fire;
  assign DispatchPlugin_logic_candidates_2_cancel = decode_ctrls_1_lane1_upIsCancel;
  assign DispatchPlugin_logic_candidates_2_ctx_valid = ((decode_ctrls_1_up_isValid && decode_ctrls_1_up_LANE_SEL_1) && (! DispatchPlugin_logic_feeds_1_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_2_ctx_laneLayerHits = {decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1,{decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1,decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1}}};
    if(decode_ctrls_1_down_TRAP_1) begin
      DispatchPlugin_logic_candidates_2_ctx_laneLayerHits = 4'b0010;
    end
  end

  assign DispatchPlugin_logic_candidates_2_ctx_uop = decode_ctrls_1_down_Decode_UOP_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY = decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER = decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH = decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 = decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 = decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 = decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_PC = decode_ctrls_1_down_PC_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_TRAP = decode_ctrls_1_down_TRAP_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID = decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE = decode_ctrls_1_down_RS1_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID = decode_ctrls_1_down_RS1_RFID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS = decode_ctrls_1_down_RS1_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE = decode_ctrls_1_down_RS2_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID = decode_ctrls_1_down_RS2_RFID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS = decode_ctrls_1_down_RS2_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE = decode_ctrls_1_down_RD_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID = decode_ctrls_1_down_RD_RFID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS = decode_ctrls_1_down_RD_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE = decode_ctrls_1_down_RS3_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID = decode_ctrls_1_down_RS3_RFID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS = decode_ctrls_1_down_RS3_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  assign when_DispatchPlugin_l368_1 = ((decode_ctrls_1_up_LANE_SEL_1 && (! DispatchPlugin_logic_feeds_1_sent)) && (! DispatchPlugin_logic_candidates_2_fire));
  assign DispatchPlugin_logic_candidates_0_ctx_valid = DispatchPlugin_logic_slots_0_ctx_valid;
  assign DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = DispatchPlugin_logic_slots_0_ctx_laneLayerHits;
  assign DispatchPlugin_logic_candidates_0_ctx_uop = DispatchPlugin_logic_slots_0_ctx_uop;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 = DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 = DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 = DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 = DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 = DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 = DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 = DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 = DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 = DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_PC = DispatchPlugin_logic_slots_0_ctx_hm_PC;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_TRAP = DispatchPlugin_logic_slots_0_ctx_hm_TRAP;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID = DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID = DispatchPlugin_logic_slots_0_ctx_hm_RS1_RFID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID = DispatchPlugin_logic_slots_0_ctx_hm_RS2_RFID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID = DispatchPlugin_logic_slots_0_ctx_hm_RD_RFID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS3_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RS3_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID = DispatchPlugin_logic_slots_0_ctx_hm_RS3_RFID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RS3_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  assign when_DispatchPlugin_l378 = (DispatchPlugin_logic_candidates_0_fire || DispatchPlugin_logic_candidates_0_cancel);
  assign _zz_GSharePlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[4 : 3];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],_zz_GSharePlugin_logic_onLearn_hash[1]} ^ _zz_GSharePlugin_logic_onLearn_hash_1);
  assign GSharePlugin_logic_onLearn_incrValue = (LearnPlugin_logic_learn_payload_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l119) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l119_1) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l119_2) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l119_3) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b00) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_onLearn_updated_1 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b01) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119_1 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1]) && (! GSharePlugin_logic_onLearn_updated_1[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1])) && GSharePlugin_logic_onLearn_updated_1[1]));
  assign GSharePlugin_logic_onLearn_updated_2 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b10) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119_2 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1]) && (! GSharePlugin_logic_onLearn_updated_2[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1])) && GSharePlugin_logic_onLearn_updated_2[1]));
  assign GSharePlugin_logic_onLearn_updated_3 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b11) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l119_3 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1]) && (! GSharePlugin_logic_onLearn_updated_3[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1])) && GSharePlugin_logic_onLearn_updated_3[1]));
  assign GSharePlugin_logic_mem_write_valid = ((LearnPlugin_logic_learn_valid && LearnPlugin_logic_learn_payload_isBranch) && (! GSharePlugin_logic_onLearn_overflow));
  assign GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
  assign GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
  assign GSharePlugin_logic_mem_write_payload_data_1 = GSharePlugin_logic_onLearn_updated_1;
  assign GSharePlugin_logic_mem_write_payload_data_2 = GSharePlugin_logic_onLearn_updated_2;
  assign GSharePlugin_logic_mem_write_payload_data_3 = GSharePlugin_logic_onLearn_updated_3;
  assign BtbPlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[21 : 10];
  always @(*) begin
    BtbPlugin_logic_memWrite_valid = (LearnPlugin_logic_learn_valid && (LearnPlugin_logic_learn_payload_badPredictedTarget && LearnPlugin_logic_learn_payload_taken));
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_valid = DecoderPlugin_logic_forgetPort_valid;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address[6:0];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address_1[6:0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_mask = (2'b01 <<< LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 2]);
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_mask = (2'b01 <<< DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[2 : 2]);
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_hash = (~ BtbPlugin_logic_onForget_hash);
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_sliceLow = LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_sliceLow = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[1 : 1];
    end
  end

  assign BtbPlugin_logic_memWrite_payload_data_0_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 1'd1);
  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPop = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_1_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_1_hash = (~ BtbPlugin_logic_onForget_hash);
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_1_sliceLow = LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_1_sliceLow = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[1 : 1];
    end
  end

  assign BtbPlugin_logic_memWrite_payload_data_1_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 1'd1);
  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_1_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_1_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_1_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_1_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_1_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_1_isPop = 1'b0;
    end
  end

  assign FpuUnpack_RS1_f32_mantissa = execute_ctrl2_up_float_RS1_lane0[22 : 0];
  assign FpuUnpack_RS1_f32_exponent = execute_ctrl2_up_float_RS1_lane0[30 : 23];
  assign FpuUnpack_RS1_f32_sign = execute_ctrl2_up_float_RS1_lane0[31];
  assign FpuUnpack_RS1_f64_mantissa = execute_ctrl2_up_float_RS1_lane0[51 : 0];
  assign FpuUnpack_RS1_f64_exponent = execute_ctrl2_up_float_RS1_lane0[62 : 52];
  assign FpuUnpack_RS1_f64_sign = execute_ctrl2_up_float_RS1_lane0[63];
  assign execute_ctrl2_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0 = (FpuUnpack_RS1_expZero && (! FpuUnpack_RS1_manZero));
  assign when_Misc_l22_9 = (execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  always @(*) begin
    if(when_Misc_l22_9) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_sign = FpuUnpack_RS1_f64_sign;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_sign = FpuUnpack_RS1_f32_sign;
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa = FpuUnpack_RS1_f64_mantissa;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa;
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS1_f64_mantissa[51];
    end else begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS1_f32_mantissa[22];
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_exponent_1;
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      FpuUnpack_RS1_manZero = (FpuUnpack_RS1_f64_mantissa == 52'h0);
    end else begin
      FpuUnpack_RS1_manZero = (FpuUnpack_RS1_f32_mantissa == 23'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      FpuUnpack_RS1_expZero = (FpuUnpack_RS1_f64_exponent == 11'h0);
    end else begin
      FpuUnpack_RS1_expZero = (FpuUnpack_RS1_f32_exponent == 8'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      FpuUnpack_RS1_expOne = (&FpuUnpack_RS1_f64_exponent);
    end else begin
      FpuUnpack_RS1_expOne = (&FpuUnpack_RS1_f32_exponent);
    end
  end

  always @(*) begin
    if(when_Misc_l22_9) begin
      FpuUnpack_RS1_recodedExpSub = 12'hc02;
    end else begin
      FpuUnpack_RS1_recodedExpSub = 12'hf82;
    end
  end

  assign switch_Misc_l245_5 = {FpuUnpack_RS1_expOne,FpuUnpack_RS1_expZero};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode = (FpuUnpack_RS1_manZero ? FloatMode_ZERO : FloatMode_NORMAL);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1 = (FpuUnpack_RS1_manZero ? FloatMode_INF : FloatMode_NAN);
  always @(*) begin
    case(switch_Misc_l245_5)
      2'b01 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_1;
      end
      default : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2 = FloatMode_NORMAL;
      end
    endcase
  end

  assign execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode_2;
  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mode;
    if(execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode = FloatMode_NAN;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_quiet;
    if(execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet = 1'b1;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_sign;
    if(execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent;
    if(FpuUnpack_RS1_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent_2;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa = execute_ctrl2_down_FpuUnpack_RS1_RS_PRE_NORM_lane0_mantissa;
    if(FpuUnpack_RS1_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa = FpuUnpack_RS1_normalizer_mantissa;
    end
  end

  assign FpuUnpack_RS1_normalizer_unpackerSel = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RS1_ENABLE_lane0) && (execute_ctrl2_down_RS1_RFID_lane0 == 1'b1)) && (! execute_ctrl2_up_TRAP_lane0));
  assign FpuUnpack_RS1_normalizer_valid = (FpuUnpack_RS1_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0);
  assign when_FpuUnpackerPlugin_l234 = (! execute_freeze_valid);
  assign when_FpuUnpackerPlugin_l235 = ((FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[0] && (! (|FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[2 : 1]))) || execute_lane0_ctrls_2_upIsCancel);
  assign when_FpuUnpackerPlugin_l236 = ((FpuUnpackerPlugin_logic_unpacker_results_0_valid && (&FpuUnpackerPlugin_logic_onUnpack_fsmServed[2 : 1])) || execute_lane0_ctrls_2_upIsCancel);
  always @(*) begin
    FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[0] = (FpuUnpack_RS1_normalizer_valid && (! FpuUnpack_RS1_normalizer_asked));
    FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[1] = (FpuUnpack_RS2_normalizer_valid && (! FpuUnpack_RS2_normalizer_asked));
    FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[2] = (FpuUnpack_RS3_normalizer_valid && (! FpuUnpack_RS3_normalizer_asked));
  end

  always @(*) begin
    FpuUnpackerPlugin_logic_onUnpack_fsmServed[0] = ((! FpuUnpack_RS1_normalizer_valid) || FpuUnpack_RS1_normalizer_served);
    FpuUnpackerPlugin_logic_onUnpack_fsmServed[1] = ((! FpuUnpack_RS2_normalizer_valid) || FpuUnpack_RS2_normalizer_served);
    FpuUnpackerPlugin_logic_onUnpack_fsmServed[2] = ((! FpuUnpack_RS3_normalizer_valid) || FpuUnpack_RS3_normalizer_served);
  end

  assign when_FpuUnpackerPlugin_l243 = FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[0];
  assign when_FpuUnpackerPlugin_l251 = (! FpuUnpack_RS1_normalizer_served);
  assign FpuUnpack_RS1_normalizer_freezeIt = ((FpuUnpack_RS1_normalizer_validReg && (! FpuUnpack_RS1_normalizer_served)) || ((FpuUnpackerPlugin_logic_onUnpack_firstCycle && FpuUnpack_RS1_normalizer_unpackerSel) && FpuUnpack_RS1_expZero));
  assign execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0 = ((execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f32_1) && (! (&execute_ctrl2_up_float_RS1_lane0[63 : 32])));
  assign FpuUnpack_RS2_f32_mantissa = execute_ctrl2_up_float_RS2_lane0[22 : 0];
  assign FpuUnpack_RS2_f32_exponent = execute_ctrl2_up_float_RS2_lane0[30 : 23];
  assign FpuUnpack_RS2_f32_sign = execute_ctrl2_up_float_RS2_lane0[31];
  assign FpuUnpack_RS2_f64_mantissa = execute_ctrl2_up_float_RS2_lane0[51 : 0];
  assign FpuUnpack_RS2_f64_exponent = execute_ctrl2_up_float_RS2_lane0[62 : 52];
  assign FpuUnpack_RS2_f64_sign = execute_ctrl2_up_float_RS2_lane0[63];
  assign execute_ctrl2_down_FpuUnpack_RS2_IS_SUBNORMAL_lane0 = (FpuUnpack_RS2_expZero && (! FpuUnpack_RS2_manZero));
  assign when_Misc_l22_10 = (execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  always @(*) begin
    if(when_Misc_l22_10) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_sign = FpuUnpack_RS2_f64_sign;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_sign = FpuUnpack_RS2_f32_sign;
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa = FpuUnpack_RS2_f64_mantissa;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa;
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS2_f64_mantissa[51];
    end else begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS2_f32_mantissa[22];
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_exponent_1;
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      FpuUnpack_RS2_manZero = (FpuUnpack_RS2_f64_mantissa == 52'h0);
    end else begin
      FpuUnpack_RS2_manZero = (FpuUnpack_RS2_f32_mantissa == 23'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      FpuUnpack_RS2_expZero = (FpuUnpack_RS2_f64_exponent == 11'h0);
    end else begin
      FpuUnpack_RS2_expZero = (FpuUnpack_RS2_f32_exponent == 8'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      FpuUnpack_RS2_expOne = (&FpuUnpack_RS2_f64_exponent);
    end else begin
      FpuUnpack_RS2_expOne = (&FpuUnpack_RS2_f32_exponent);
    end
  end

  always @(*) begin
    if(when_Misc_l22_10) begin
      FpuUnpack_RS2_recodedExpSub = 12'hc02;
    end else begin
      FpuUnpack_RS2_recodedExpSub = 12'hf82;
    end
  end

  assign switch_Misc_l245_6 = {FpuUnpack_RS2_expOne,FpuUnpack_RS2_expZero};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode = (FpuUnpack_RS2_manZero ? FloatMode_ZERO : FloatMode_NORMAL);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1 = (FpuUnpack_RS2_manZero ? FloatMode_INF : FloatMode_NAN);
  always @(*) begin
    case(switch_Misc_l245_6)
      2'b01 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_1;
      end
      default : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2 = FloatMode_NORMAL;
      end
    endcase
  end

  assign execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode_2;
  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mode;
    if(execute_ctrl2_down_FpuUnpack_RS2_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode = FloatMode_NAN;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_quiet;
    if(execute_ctrl2_down_FpuUnpack_RS2_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet = 1'b1;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_sign;
    if(execute_ctrl2_down_FpuUnpack_RS2_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent;
    if(FpuUnpack_RS2_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_exponent_2;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa = execute_ctrl2_down_FpuUnpack_RS2_RS_PRE_NORM_lane0_mantissa;
    if(FpuUnpack_RS2_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa = FpuUnpack_RS2_normalizer_mantissa;
    end
  end

  assign FpuUnpack_RS2_normalizer_unpackerSel = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RS2_ENABLE_lane0) && (execute_ctrl2_down_RS2_RFID_lane0 == 1'b1)) && (! execute_ctrl2_up_TRAP_lane0));
  assign FpuUnpack_RS2_normalizer_valid = (FpuUnpack_RS2_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS2_IS_SUBNORMAL_lane0);
  assign when_FpuUnpackerPlugin_l234_1 = (! execute_freeze_valid);
  assign when_FpuUnpackerPlugin_l235_1 = ((FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[1] && (! (|FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[2 : 2]))) || execute_lane0_ctrls_2_upIsCancel);
  assign when_FpuUnpackerPlugin_l236_1 = ((FpuUnpackerPlugin_logic_unpacker_results_0_valid && (&FpuUnpackerPlugin_logic_onUnpack_fsmServed[2 : 2])) || execute_lane0_ctrls_2_upIsCancel);
  assign when_FpuUnpackerPlugin_l243_1 = FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[1];
  assign when_FpuUnpackerPlugin_l251_1 = (! FpuUnpack_RS2_normalizer_served);
  assign FpuUnpack_RS2_normalizer_freezeIt = ((FpuUnpack_RS2_normalizer_validReg && (! FpuUnpack_RS2_normalizer_served)) || ((FpuUnpackerPlugin_logic_onUnpack_firstCycle && FpuUnpack_RS2_normalizer_unpackerSel) && FpuUnpack_RS2_expZero));
  assign execute_ctrl2_down_FpuUnpack_RS2_badBoxing_HIT_lane0 = ((execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f32_1) && (! (&execute_ctrl2_up_float_RS2_lane0[63 : 32])));
  assign FpuUnpack_RS3_f32_mantissa = execute_ctrl2_up_float_RS3_lane0[22 : 0];
  assign FpuUnpack_RS3_f32_exponent = execute_ctrl2_up_float_RS3_lane0[30 : 23];
  assign FpuUnpack_RS3_f32_sign = execute_ctrl2_up_float_RS3_lane0[31];
  assign FpuUnpack_RS3_f64_mantissa = execute_ctrl2_up_float_RS3_lane0[51 : 0];
  assign FpuUnpack_RS3_f64_exponent = execute_ctrl2_up_float_RS3_lane0[62 : 52];
  assign FpuUnpack_RS3_f64_sign = execute_ctrl2_up_float_RS3_lane0[63];
  assign execute_ctrl2_down_FpuUnpack_RS3_IS_SUBNORMAL_lane0 = (FpuUnpack_RS3_expZero && (! FpuUnpack_RS3_manZero));
  assign when_Misc_l22_11 = (execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  always @(*) begin
    if(when_Misc_l22_11) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_sign = FpuUnpack_RS3_f64_sign;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_sign = FpuUnpack_RS3_f32_sign;
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa = FpuUnpack_RS3_f64_mantissa;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa;
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS3_f64_mantissa[51];
    end else begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_quiet = FpuUnpack_RS3_f32_mantissa[22];
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent;
    end else begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_exponent_1;
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      FpuUnpack_RS3_manZero = (FpuUnpack_RS3_f64_mantissa == 52'h0);
    end else begin
      FpuUnpack_RS3_manZero = (FpuUnpack_RS3_f32_mantissa == 23'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      FpuUnpack_RS3_expZero = (FpuUnpack_RS3_f64_exponent == 11'h0);
    end else begin
      FpuUnpack_RS3_expZero = (FpuUnpack_RS3_f32_exponent == 8'h0);
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      FpuUnpack_RS3_expOne = (&FpuUnpack_RS3_f64_exponent);
    end else begin
      FpuUnpack_RS3_expOne = (&FpuUnpack_RS3_f32_exponent);
    end
  end

  always @(*) begin
    if(when_Misc_l22_11) begin
      FpuUnpack_RS3_recodedExpSub = 12'hc02;
    end else begin
      FpuUnpack_RS3_recodedExpSub = 12'hf82;
    end
  end

  assign switch_Misc_l245_7 = {FpuUnpack_RS3_expOne,FpuUnpack_RS3_expZero};
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode = (FpuUnpack_RS3_manZero ? FloatMode_ZERO : FloatMode_NORMAL);
  assign _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1 = (FpuUnpack_RS3_manZero ? FloatMode_INF : FloatMode_NAN);
  always @(*) begin
    case(switch_Misc_l245_7)
      2'b01 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2 = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_1;
      end
      default : begin
        _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2 = FloatMode_NORMAL;
      end
    endcase
  end

  assign execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode_2;
  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mode;
    if(execute_ctrl2_down_FpuUnpack_RS3_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode = FloatMode_NAN;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_quiet = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_quiet;
    if(execute_ctrl2_down_FpuUnpack_RS3_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_quiet = 1'b1;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_sign = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_sign;
    if(execute_ctrl2_down_FpuUnpack_RS3_badBoxing_HIT_lane0) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_sign = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent;
    if(FpuUnpack_RS3_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent = _zz_execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_exponent_2;
    end
  end

  always @(*) begin
    execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mantissa = execute_ctrl2_down_FpuUnpack_RS3_RS_PRE_NORM_lane0_mantissa;
    if(FpuUnpack_RS3_normalizer_asked) begin
      execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mantissa = FpuUnpack_RS3_normalizer_mantissa;
    end
  end

  assign FpuUnpack_RS3_normalizer_unpackerSel = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RS3_ENABLE_lane0) && (execute_ctrl2_down_RS3_RFID_lane0 == 1'b1)) && (! execute_ctrl2_up_TRAP_lane0));
  assign FpuUnpack_RS3_normalizer_valid = (FpuUnpack_RS3_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS3_IS_SUBNORMAL_lane0);
  assign when_FpuUnpackerPlugin_l234_2 = (! execute_freeze_valid);
  assign when_FpuUnpackerPlugin_l235_2 = ((FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[2] && (! 1'b0)) || execute_lane0_ctrls_2_upIsCancel);
  assign when_FpuUnpackerPlugin_l236_2 = ((FpuUnpackerPlugin_logic_unpacker_results_0_valid && 1'b1) || execute_lane0_ctrls_2_upIsCancel);
  assign when_FpuUnpackerPlugin_l243_2 = FpuUnpackerPlugin_logic_onUnpack_fsmRequesters[2];
  assign when_FpuUnpackerPlugin_l251_2 = (! FpuUnpack_RS3_normalizer_served);
  assign FpuUnpack_RS3_normalizer_freezeIt = ((FpuUnpack_RS3_normalizer_validReg && (! FpuUnpack_RS3_normalizer_served)) || ((FpuUnpackerPlugin_logic_onUnpack_firstCycle && FpuUnpack_RS3_normalizer_unpackerSel) && FpuUnpack_RS3_expZero));
  assign execute_ctrl2_down_FpuUnpack_RS3_badBoxing_HIT_lane0 = ((execute_ctrl2_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f32_1) && (! (&execute_ctrl2_up_float_RS3_lane0[63 : 32])));
  assign FpuUnpackerPlugin_logic_unpackDone = (! (|{FpuUnpack_RS3_normalizer_freezeIt,{FpuUnpack_RS2_normalizer_freezeIt,FpuUnpack_RS1_normalizer_freezeIt}}));
  assign FpuUnpackerPlugin_logic_onCvt_rs1Zero = (execute_ctrl2_up_integer_RS1_lane0[31 : 0] == 32'h0);
  assign FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_valid = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuUnpackerPlugin_SEL_I2F_lane0) && FpuUnpackerPlugin_logic_unpackDone) && (! FpuUnpackerPlugin_logic_onCvt_asked));
  assign FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_payload_data = {20'd0, _zz_io_inputs_1_payload_data};
  assign FpuUnpackerPlugin_logic_onCvt_freezeIt = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuUnpackerPlugin_SEL_I2F_lane0) && (! FpuUnpackerPlugin_logic_onCvt_served));
  assign FpuUnpackerPlugin_logic_packPort_cmd_at[0] = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuUnpackerPlugin_SEL_I2F_lane0);
  assign _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX = 5'h0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_flags_NX = _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX[0];
  assign FpuUnpackerPlugin_logic_packPort_cmd_flags_UF = _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX[1];
  assign FpuUnpackerPlugin_logic_packPort_cmd_flags_OF = _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX[2];
  assign FpuUnpackerPlugin_logic_packPort_cmd_flags_DZ = _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX[3];
  assign FpuUnpackerPlugin_logic_packPort_cmd_flags_NV = _zz_FpuUnpackerPlugin_logic_packPort_cmd_flags_NX[4];
  assign FpuUnpackerPlugin_logic_packPort_cmd_format = execute_ctrl2_down_FpuUtils_FORMAT_lane0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_roundMode = execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_value_quiet = 1'b0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_value_sign = execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  assign FpuUnpackerPlugin_logic_packPort_cmd_value_exponent = _zz_FpuUnpackerPlugin_logic_packPort_cmd_value_exponent;
  assign FpuUnpackerPlugin_logic_packPort_cmd_value_mantissa = ({2'd0,FpuUnpackerPlugin_logic_onCvt_fsmResult_data} <<< 2'd2);
  always @(*) begin
    FpuUnpackerPlugin_logic_packPort_cmd_value_mode = FloatMode_NORMAL;
    if(FpuUnpackerPlugin_logic_onCvt_rs1Zero) begin
      FpuUnpackerPlugin_logic_packPort_cmd_value_mode = FloatMode_ZERO;
    end
  end

  assign FpuUnpackerPlugin_logic_unpacker_node_0_isValid = FpuUnpackerPlugin_logic_unpacker_node_0_valid;
  assign FpuUnpackerPlugin_logic_unpacker_node_1_isValid = FpuUnpackerPlugin_logic_unpacker_node_1_valid;
  assign FpuUnpackerPlugin_logic_unpacker_node_2_isValid = FpuUnpackerPlugin_logic_unpacker_node_2_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_hits = {lane0_IntFormatPlugin_logic_stages_0_wb_valid,early0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early0_BranchPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane0_IntFormatPlugin_logic_stages_0_wb_payload : 32'h0));
  assign execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_0_hits)) && execute_ctrl2_up_RD_ENABLE_lane0) && execute_ctrl2_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_hits = lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_muxed = (lane0_integer_WriteBackPlugin_logic_stages_1_hits[0] ? lane0_IntFormatPlugin_logic_stages_2_wb_payload : 32'h0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_merged = (execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_1_hits)) && execute_ctrl3_up_RD_ENABLE_lane0) && execute_ctrl3_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_hits = {lane0_IntFormatPlugin_logic_stages_1_wb_valid,late0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_2_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_2_hits[0] ? late0_BranchPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_2_hits[1] ? lane0_IntFormatPlugin_logic_stages_1_wb_payload : 32'h0));
  assign lane0_integer_WriteBackPlugin_logic_stages_2_merged = (execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_2_muxed);
  assign execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_valid = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_2_hits)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  assign lane0_integer_WriteBackPlugin_logic_write_port_valid = (((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_write_port_address = execute_ctrl4_down_RD_PHYS_lane0[4 : 0];
  assign lane0_integer_WriteBackPlugin_logic_write_port_data = execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_hits = {lane1_IntFormatPlugin_logic_stages_0_wb_valid,early1_BranchPlugin_logic_wb_valid};
  assign lane1_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane1_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early1_BranchPlugin_logic_wb_payload : 32'h0) | (lane1_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane1_IntFormatPlugin_logic_stages_0_wb_payload : 32'h0));
  assign execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass = lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((execute_ctrl2_down_LANE_SEL_lane1 && execute_ctrl2_down_isReady) && (! execute_lane1_ctrls_2_downIsCancel)) && (|lane1_integer_WriteBackPlugin_logic_stages_0_hits)) && execute_ctrl2_up_RD_ENABLE_lane1) && execute_ctrl2_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_hits = {lane1_IntFormatPlugin_logic_stages_1_wb_valid,late1_BranchPlugin_logic_wb_valid};
  assign lane1_integer_WriteBackPlugin_logic_stages_1_muxed = ((lane1_integer_WriteBackPlugin_logic_stages_1_hits[0] ? late1_BranchPlugin_logic_wb_payload : 32'h0) | (lane1_integer_WriteBackPlugin_logic_stages_1_hits[1] ? lane1_IntFormatPlugin_logic_stages_1_wb_payload : 32'h0));
  assign lane1_integer_WriteBackPlugin_logic_stages_1_merged = (execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 | lane1_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass = lane1_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((execute_ctrl4_down_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_downIsCancel)) && (|lane1_integer_WriteBackPlugin_logic_stages_1_hits)) && execute_ctrl4_up_RD_ENABLE_lane1) && execute_ctrl4_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane1_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane1_integer_WriteBackPlugin_logic_write_port_valid = (((((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_upIsCancel)) && execute_ctrl4_up_RD_ENABLE_lane1) && execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1) && execute_ctrl4_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_write_port_address = execute_ctrl4_down_RD_PHYS_lane1[4 : 0];
  assign lane1_integer_WriteBackPlugin_logic_write_port_data = execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  assign lane1_integer_WriteBackPlugin_logic_write_port_uopId = execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign lane0_float_WriteBackPlugin_logic_stages_0_hits = FpuCmpPlugin_logic_fwb_valid;
  assign lane0_float_WriteBackPlugin_logic_stages_0_muxed = (lane0_float_WriteBackPlugin_logic_stages_0_hits[0] ? FpuCmpPlugin_logic_fwb_payload : 64'h0);
  assign execute_ctrl3_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_0_write_valid = (((((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_0_hits)) && execute_ctrl3_up_RD_ENABLE_lane0) && execute_ctrl3_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_0_write_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_0_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_1_hits = {FpuPackerPlugin_wb_at_2_valid,{FpuMvPlugin_logic_fwb_valid,LsuPlugin_logic_fpwb_valid}};
  assign lane0_float_WriteBackPlugin_logic_stages_1_muxed = (((lane0_float_WriteBackPlugin_logic_stages_1_hits[0] ? LsuPlugin_logic_fpwb_payload : 64'h0) | (lane0_float_WriteBackPlugin_logic_stages_1_hits[1] ? FpuMvPlugin_logic_fwb_payload : 64'h0)) | (lane0_float_WriteBackPlugin_logic_stages_1_hits[2] ? FpuPackerPlugin_wb_at_2_payload : 64'h0));
  assign lane0_float_WriteBackPlugin_logic_stages_1_merged = (execute_ctrl4_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 | lane0_float_WriteBackPlugin_logic_stages_1_muxed);
  assign execute_ctrl4_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_1_merged;
  assign lane0_float_WriteBackPlugin_logic_stages_1_write_valid = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_1_hits)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_1_write_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_1_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_1_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_2_hits = FpuPackerPlugin_wb_at_3_valid;
  assign lane0_float_WriteBackPlugin_logic_stages_2_muxed = (lane0_float_WriteBackPlugin_logic_stages_2_hits[0] ? FpuPackerPlugin_wb_at_3_payload : 64'h0);
  assign lane0_float_WriteBackPlugin_logic_stages_2_merged = (execute_ctrl5_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 | lane0_float_WriteBackPlugin_logic_stages_2_muxed);
  assign execute_ctrl5_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_2_merged;
  assign lane0_float_WriteBackPlugin_logic_stages_2_write_valid = (((((execute_ctrl5_down_LANE_SEL_lane0 && execute_ctrl5_down_isReady) && (! execute_lane0_ctrls_5_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_2_hits)) && execute_ctrl5_up_RD_ENABLE_lane0) && execute_ctrl5_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_2_write_payload_uopId = execute_ctrl5_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_2_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_2_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_3_hits = FpuPackerPlugin_wb_at_5_valid;
  assign lane0_float_WriteBackPlugin_logic_stages_3_muxed = (lane0_float_WriteBackPlugin_logic_stages_3_hits[0] ? FpuPackerPlugin_wb_at_5_payload : 64'h0);
  assign lane0_float_WriteBackPlugin_logic_stages_3_merged = (execute_ctrl7_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 | lane0_float_WriteBackPlugin_logic_stages_3_muxed);
  assign execute_ctrl7_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_3_merged;
  assign lane0_float_WriteBackPlugin_logic_stages_3_write_valid = (((((execute_ctrl7_down_LANE_SEL_lane0 && execute_ctrl7_down_isReady) && (! execute_lane0_ctrls_7_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_3_hits)) && execute_ctrl7_up_RD_ENABLE_lane0) && execute_ctrl7_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_3_write_payload_uopId = execute_ctrl7_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_3_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_3_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_4_hits = FpuPackerPlugin_wb_at_6_valid;
  assign lane0_float_WriteBackPlugin_logic_stages_4_muxed = (lane0_float_WriteBackPlugin_logic_stages_4_hits[0] ? FpuPackerPlugin_wb_at_6_payload : 64'h0);
  assign lane0_float_WriteBackPlugin_logic_stages_4_merged = (execute_ctrl8_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 | lane0_float_WriteBackPlugin_logic_stages_4_muxed);
  assign execute_ctrl8_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_4_merged;
  assign lane0_float_WriteBackPlugin_logic_stages_4_write_valid = (((((execute_ctrl8_down_LANE_SEL_lane0 && execute_ctrl8_down_isReady) && (! execute_lane0_ctrls_8_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_4_hits)) && execute_ctrl8_up_RD_ENABLE_lane0) && execute_ctrl8_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_4_write_payload_uopId = execute_ctrl8_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_4_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_4_muxed;
  assign lane0_float_WriteBackPlugin_logic_stages_5_hits = FpuPackerPlugin_wb_at_9_valid;
  assign lane0_float_WriteBackPlugin_logic_stages_5_muxed = (lane0_float_WriteBackPlugin_logic_stages_5_hits[0] ? FpuPackerPlugin_wb_at_9_payload : 64'h0);
  assign lane0_float_WriteBackPlugin_logic_stages_5_merged = (execute_ctrl11_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 | lane0_float_WriteBackPlugin_logic_stages_5_muxed);
  assign execute_ctrl11_lane0_float_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_float_WriteBackPlugin_logic_stages_5_merged;
  assign lane0_float_WriteBackPlugin_logic_stages_5_write_valid = (((((execute_ctrl11_down_LANE_SEL_lane0 && execute_ctrl11_down_isReady) && (! execute_lane0_ctrls_11_downIsCancel)) && (|lane0_float_WriteBackPlugin_logic_stages_5_hits)) && execute_ctrl11_up_RD_ENABLE_lane0) && execute_ctrl11_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_stages_5_write_payload_uopId = execute_ctrl11_down_Decode_UOP_ID_lane0;
  assign lane0_float_WriteBackPlugin_logic_stages_5_write_payload_data = lane0_float_WriteBackPlugin_logic_stages_5_muxed;
  assign lane0_float_WriteBackPlugin_logic_write_port_valid = (((((execute_ctrl11_up_LANE_SEL_lane0 && execute_ctrl11_down_isReady) && (! execute_lane0_ctrls_11_upIsCancel)) && execute_ctrl11_up_RD_ENABLE_lane0) && execute_ctrl11_down_lane0_float_WriteBackPlugin_SEL_lane0) && execute_ctrl11_down_COMMIT_lane0);
  assign lane0_float_WriteBackPlugin_logic_write_port_address = execute_ctrl11_down_RD_PHYS_lane0[4 : 0];
  assign lane0_float_WriteBackPlugin_logic_write_port_data = execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  assign lane0_float_WriteBackPlugin_logic_write_port_uopId = execute_ctrl11_down_Decode_UOP_ID_lane0;
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00003064) == 32'h00003000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00106060) == 32'h00006000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h000060e0) == 32'h00006080);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006860) == 32'h00006800);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006160) == 32'h00006100);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00406060) == 32'h00406000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_7 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006260) == 32'h00006200);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_8 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h01006060) == 32'h01006000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00806060) == 32'h00806000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006460) == 32'h00006400);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_11 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002070) == 32'h00000010);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_12 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00004070) == 32'h00000010);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_13 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h02000070) == 32'h00000030);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_14 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000074) == 32'h00000060);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000068) == 32'h00000068);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_16[0];
  assign decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002070) == 32'h00002070);
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001070) == 32'h00001070);
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h70000070) == 32'h00000050);
  assign decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_0[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_0_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_0[0];
  assign decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_0[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_0_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_0[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00003064) == 32'h00003000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00106060) == 32'h00006000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h000060e0) == 32'h00006080);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006860) == 32'h00006800);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006160) == 32'h00006100);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00406060) == 32'h00406000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_7 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006260) == 32'h00006200);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_8 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h01006060) == 32'h01006000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00806060) == 32'h00806000);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006460) == 32'h00006400);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_11 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002070) == 32'h00000010);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_12 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00004070) == 32'h00000010);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_13 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h02000070) == 32'h00000030);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_14 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000074) == 32'h00000060);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000068) == 32'h00000068);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_16[0];
  assign decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002070) == 32'h00002070);
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001070) == 32'h00001070);
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1[0];
  assign _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h70000070) == 32'h00000050);
  assign decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_1_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_1[0];
  assign decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1 = _zz_decode_ctrls_1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_1_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_2_1[0];
  assign decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1 = _zz_decode_ctrls_1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_1[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1[0];
  always @(*) begin
    FpuClassPlugin_logic_onWb_fclassResult = 10'h0;
    FpuClassPlugin_logic_onWb_fclassResult[0] = (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF));
    FpuClassPlugin_logic_onWb_fclassResult[1] = ((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NORMAL)) && (! execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0));
    FpuClassPlugin_logic_onWb_fclassResult[2] = ((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NORMAL)) && execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0);
    FpuClassPlugin_logic_onWb_fclassResult[3] = (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO));
    FpuClassPlugin_logic_onWb_fclassResult[4] = ((! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign) && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO));
    FpuClassPlugin_logic_onWb_fclassResult[5] = (((! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign) && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NORMAL)) && execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0);
    FpuClassPlugin_logic_onWb_fclassResult[6] = (((! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign) && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NORMAL)) && (! execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0));
    FpuClassPlugin_logic_onWb_fclassResult[7] = ((! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign) && (execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF));
    FpuClassPlugin_logic_onWb_fclassResult[8] = ((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet));
    FpuClassPlugin_logic_onWb_fclassResult[9] = ((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet);
  end

  assign FpuClassPlugin_logic_onWb_expSubnormal = ((execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1) ? 11'h401 : 11'h781);
  assign FpuClassPlugin_logic_iwb_valid = execute_ctrl3_down_FpuClassPlugin_SEL_lane0;
  assign FpuClassPlugin_logic_iwb_payload = {22'd0, FpuClassPlugin_logic_onWb_fclassResult};
  assign FpuCmpPlugin_logic_onCmp_signalQuiet = (execute_ctrl2_down_FpuCmpPlugin_SEL_CMP_lane0 && execute_ctrl2_down_FpuCmpPlugin_LESS_lane0);
  assign FpuCmpPlugin_logic_onCmp_rs1NanNv = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && ((! execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet) || FpuCmpPlugin_logic_onCmp_signalQuiet));
  assign FpuCmpPlugin_logic_onCmp_rs2NanNv = ((execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN) && ((! execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet) || FpuCmpPlugin_logic_onCmp_signalQuiet));
  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_NV_lane0 = (FpuCmpPlugin_logic_onCmp_rs1NanNv || FpuCmpPlugin_logic_onCmp_rs2NanNv);
  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_bothZero_lane0 = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO) && (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO));
  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0 = ($signed(_zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0) == $signed(_zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0_1));
  always @(*) begin
    execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1Equal_lane0 = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign == execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign) && execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0) && (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa == execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa));
    if(when_FpuCmpPlugin_l114) begin
      execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1Equal_lane0 = 1'b1;
    end
  end

  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0 = ($signed(_zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0) < $signed(_zz_execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0_1));
  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1MantissaSmaller_lane0 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa < execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa);
  always @(*) begin
    FpuCmpPlugin_logic_onCmp_rs1AbsSmaller = (execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1ExpSmaller_lane0 || (execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_expEqual_lane0 && execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1MantissaSmaller_lane0));
    if(when_FpuCmpPlugin_l110) begin
      FpuCmpPlugin_logic_onCmp_rs1AbsSmaller = 1'b1;
    end
    if(when_FpuCmpPlugin_l111) begin
      FpuCmpPlugin_logic_onCmp_rs1AbsSmaller = 1'b1;
    end
    if(when_FpuCmpPlugin_l112) begin
      FpuCmpPlugin_logic_onCmp_rs1AbsSmaller = 1'b0;
    end
    if(when_FpuCmpPlugin_l113) begin
      FpuCmpPlugin_logic_onCmp_rs1AbsSmaller = 1'b0;
    end
  end

  assign when_FpuCmpPlugin_l110 = (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF);
  assign when_FpuCmpPlugin_l111 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO);
  assign when_FpuCmpPlugin_l112 = (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO);
  assign when_FpuCmpPlugin_l113 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF);
  assign when_FpuCmpPlugin_l114 = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign == execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign) && (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF)) && (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF));
  assign switch_Misc_l245_8 = {execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign,execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign};
  always @(*) begin
    case(switch_Misc_l245_8)
      2'b00 : begin
        FpuCmpPlugin_logic_onCmp_rs1Smaller = FpuCmpPlugin_logic_onCmp_rs1AbsSmaller;
      end
      2'b01 : begin
        FpuCmpPlugin_logic_onCmp_rs1Smaller = 1'b0;
      end
      2'b10 : begin
        FpuCmpPlugin_logic_onCmp_rs1Smaller = 1'b1;
      end
      default : begin
        FpuCmpPlugin_logic_onCmp_rs1Smaller = ((! FpuCmpPlugin_logic_onCmp_rs1AbsSmaller) && (! execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1Equal_lane0));
      end
    endcase
  end

  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0 = (! (((FpuCmpPlugin_logic_onCmp_rs1Smaller ^ (! execute_ctrl2_down_FpuCmpPlugin_LESS_lane0)) && (! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN))) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN)));
  always @(*) begin
    execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0 = (((FpuCmpPlugin_logic_onCmp_rs1Smaller && (! execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_bothZero_lane0)) && execute_ctrl2_down_FpuCmpPlugin_LESS_lane0) || ((execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_rs1Equal_lane0 || execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_bothZero_lane0) && execute_ctrl2_down_FpuCmpPlugin_EQUAL_lane0));
    if(when_FpuCmpPlugin_l124) begin
      execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0 = 1'b0;
    end
  end

  assign when_FpuCmpPlugin_l124 = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN));
  assign execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0 = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign && execute_ctrl2_down_FpuCmpPlugin_SGNJ_RS1_lane0) ^ execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign) ^ execute_ctrl2_down_FpuCmpPlugin_INVERT_lane0);
  assign FpuCmpPlugin_logic_ffwb_ats[0] = ((execute_ctrl2_down_FpuCmpPlugin_SEL_FLOAT_lane0 && (execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0 == FpuCmpFloatOp_MIN_MAX)) || execute_ctrl2_down_FpuCmpPlugin_SEL_CMP_lane0);
  assign FpuCmpPlugin_logic_ffwb_flags_NX = 1'b0;
  assign FpuCmpPlugin_logic_ffwb_flags_UF = 1'b0;
  assign FpuCmpPlugin_logic_ffwb_flags_OF = 1'b0;
  assign FpuCmpPlugin_logic_ffwb_flags_DZ = 1'b0;
  assign FpuCmpPlugin_logic_ffwb_flags_NV = execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_NV_lane0;
  assign FpuCmpPlugin_logic_iwb_valid = execute_ctrl3_down_FpuCmpPlugin_SEL_CMP_lane0;
  assign FpuCmpPlugin_logic_iwb_payload = {31'd0, _zz_FpuCmpPlugin_logic_iwb_payload};
  assign FpuCmpPlugin_logic_fwb_valid = execute_ctrl3_down_FpuCmpPlugin_SEL_FLOAT_lane0;
  always @(*) begin
    FpuCmpPlugin_logic_fwb_payload = (((execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0 == FpuCmpFloatOp_MIN_MAX) && execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0) ? execute_ctrl3_up_float_RS2_lane0 : execute_ctrl3_up_float_RS1_lane0);
    if(FpuCmpPlugin_logic_onFloatWb_doNan) begin
      if(when_Misc_l22_12) begin
        FpuCmpPlugin_logic_fwb_payload[62 : 52] = 11'h7ff;
      end else begin
        FpuCmpPlugin_logic_fwb_payload[30 : 23] = 8'hff;
      end
      if(when_Misc_l22_13) begin
        FpuCmpPlugin_logic_fwb_payload[51 : 0] = 52'h0;
      end else begin
        FpuCmpPlugin_logic_fwb_payload[22 : 0] = 23'h0;
      end
      if(when_Misc_l22_14) begin
        FpuCmpPlugin_logic_fwb_payload[51] = 1'b1;
      end else begin
        FpuCmpPlugin_logic_fwb_payload[22] = 1'b1;
      end
      if(when_Misc_l22_15) begin
        FpuCmpPlugin_logic_fwb_payload[63] = 1'b0;
      end else begin
        FpuCmpPlugin_logic_fwb_payload[31] = 1'b0;
      end
      if(when_FpuCmpPlugin_l149) begin
        FpuCmpPlugin_logic_fwb_payload[63 : 32] = 32'hffffffff;
      end
    end
    if(when_FpuCmpPlugin_l153) begin
      if(when_Misc_l22_16) begin
        FpuCmpPlugin_logic_fwb_payload[63] = execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
      end else begin
        FpuCmpPlugin_logic_fwb_payload[31] = execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
      end
    end
  end

  always @(*) begin
    FpuCmpPlugin_logic_onFloatWb_doNan = (((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN)) && (execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0 == FpuCmpFloatOp_MIN_MAX));
    if(when_FpuCmpPlugin_l153) begin
      if(execute_ctrl3_down_FpuUnpack_RS1_badBoxing_HIT_lane0) begin
        FpuCmpPlugin_logic_onFloatWb_doNan = 1'b1;
      end
    end
  end

  assign when_Misc_l22_12 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_13 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_14 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_Misc_l22_15 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign when_FpuCmpPlugin_l149 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f32_1);
  assign when_FpuCmpPlugin_l153 = (execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0 == FpuCmpFloatOp_SGNJ);
  assign when_Misc_l22_16 = (execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f64_1);
  assign execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0 = _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0;
  assign _zz_when_UInt_l119 = execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShiftFull_lane0;
  assign when_UInt_l119_3 = (|_zz_when_UInt_l119[11 : 6]);
  always @(*) begin
    if(when_UInt_l119_3) begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 = 6'h3f;
    end else begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 = _zz_when_UInt_l119[5 : 0];
    end
  end

  assign execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 = _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  assign _zz_when_Utils_l1585_16 = {{1'b1,execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa},1'b0};
  assign _zz_when_Utils_l1585_17 = execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0[3 : 0];
  always @(*) begin
    _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = 1'b0;
    if(when_Utils_l1585_13) begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = 1'b1;
    end
    if(when_Utils_l1585_14) begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = 1'b1;
    end
    if(when_Utils_l1585_15) begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = 1'b1;
    end
    if(when_Utils_l1585_16) begin
      _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1 = 1'b1;
    end
  end

  assign when_Utils_l1585_13 = (_zz_when_Utils_l1585_17[0] && (_zz_when_Utils_l1585_16[0 : 0] != 1'b0));
  assign when_Utils_l1585_14 = (_zz_when_Utils_l1585_17[1] && (_zz_when_Utils_l1585_2[1 : 0] != 2'b00));
  assign when_Utils_l1585_15 = (_zz_when_Utils_l1585_17[2] && (_zz_when_Utils_l1585_1[3 : 0] != 4'b0000));
  assign when_Utils_l1585_16 = (_zz_when_Utils_l1585_17[3] && (_zz_when_Utils_l1585[7 : 0] != 8'h0));
  assign execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 = (_zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 | _zz_execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2);
  assign FpuF2iPlugin_logic_onShift_signed = (! execute_ctrl3_down_Decode_UOP_lane0[20]);
  assign _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6 = ({4'd0,_zz__zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6} <<< 3'd4);
  always @(*) begin
    _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b0;
    if(when_Utils_l1585_17) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
    if(when_Utils_l1585_18) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
    if(when_Utils_l1585_19) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
    if(when_Utils_l1585_20) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
    if(when_Utils_l1585_21) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
    if(when_Utils_l1585_22) begin
      _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = 1'b1;
    end
  end

  assign when_Utils_l1585_17 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[0] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0[0 : 0] != 1'b0));
  assign when_Utils_l1585_18 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[1] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_1[1 : 0] != 2'b00));
  assign when_Utils_l1585_19 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[2] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_2[3 : 0] != 4'b0000));
  assign when_Utils_l1585_20 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[3] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_3[7 : 0] != 8'h0));
  assign when_Utils_l1585_21 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[4] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_4[15 : 0] != 16'h0));
  assign when_Utils_l1585_22 = (_zz_execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6[5] && (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_5[31 : 0] != 32'h0));
  assign execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = (execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0_6 | _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0_1);
  assign FpuF2iPlugin_logic_onShift_high = execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0[53 : 22];
  assign FpuF2iPlugin_logic_onShift_low = execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0[21 : 0];
  assign FpuF2iPlugin_logic_onShift_unsigned = FpuF2iPlugin_logic_onShift_high;
  assign FpuF2iPlugin_logic_onShift_round = {FpuF2iPlugin_logic_onShift_low[21],(|FpuF2iPlugin_logic_onShift_low[20 : 0])};
  assign execute_ctrl3_down_FpuF2iPlugin_logic_onShift_resign_lane0 = (FpuF2iPlugin_logic_onShift_signed && execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign);
  always @(*) begin
    case(execute_ctrl3_down_FpuUtils_ROUNDING_lane0)
      FpuRoundMode_RNE : begin
        _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = (FpuF2iPlugin_logic_onShift_round[1] && (FpuF2iPlugin_logic_onShift_round[0] || FpuF2iPlugin_logic_onShift_unsigned[0]));
      end
      FpuRoundMode_RTZ : begin
        _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = 1'b0;
      end
      FpuRoundMode_RDN : begin
        _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = ((FpuF2iPlugin_logic_onShift_round != 2'b00) && execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign);
      end
      FpuRoundMode_RUP : begin
        _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = ((FpuF2iPlugin_logic_onShift_round != 2'b00) && (! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign));
      end
      default : begin
        _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = FpuF2iPlugin_logic_onShift_round[1];
      end
    endcase
  end

  assign execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0 = _zz_execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0;
  assign execute_ctrl3_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0 = (execute_ctrl3_down_FpuF2iPlugin_logic_onShift_resign_lane0 ^ execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0);
  assign FpuF2iPlugin_logic_onResult_signed = (! execute_ctrl4_down_Decode_UOP_lane0[20]);
  assign FpuF2iPlugin_logic_onResult_i64 = execute_ctrl4_down_Decode_UOP_lane0[21];
  assign FpuF2iPlugin_logic_onResult_high = execute_ctrl4_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0[53 : 22];
  assign FpuF2iPlugin_logic_onResult_low = execute_ctrl4_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0[21 : 0];
  assign FpuF2iPlugin_logic_onResult_unsigned = FpuF2iPlugin_logic_onResult_high;
  assign FpuF2iPlugin_logic_onResult_round = {FpuF2iPlugin_logic_onResult_low[21],(|FpuF2iPlugin_logic_onResult_low[20 : 0])};
  assign FpuF2iPlugin_logic_onResult_halfRater_freezeIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_FpuF2iPlugin_SEL_lane0) && FpuF2iPlugin_logic_onResult_halfRater_firstCycle);
  always @(*) begin
    FpuF2iPlugin_logic_onResult_resultRaw = FpuF2iPlugin_logic_onResult_inverter;
    if(FpuF2iPlugin_logic_onResult_isZero) begin
      FpuF2iPlugin_logic_onResult_resultRaw = 32'h0;
    end else begin
      if(when_FpuF2iPlugin_l129) begin
        FpuF2iPlugin_logic_onResult_resultRaw = (FpuF2iPlugin_logic_onResult_overflow ? 32'hffffffff : 32'h0);
        FpuF2iPlugin_logic_onResult_resultRaw[31] = (FpuF2iPlugin_logic_onResult_signed ^ FpuF2iPlugin_logic_onResult_overflow);
      end
    end
  end

  assign _zz_FpuF2iPlugin_logic_onResult_expMax[0] = (! FpuF2iPlugin_logic_onResult_signed);
  assign FpuF2iPlugin_logic_onResult_expMax = _zz_FpuF2iPlugin_logic_onResult_expMax_1;
  assign FpuF2iPlugin_logic_onResult_expMin = (FpuF2iPlugin_logic_onResult_i64 ? 6'h3f : _zz_FpuF2iPlugin_logic_onResult_expMin);
  assign FpuF2iPlugin_logic_onResult_unsignedMin = 32'h80000000;
  always @(*) begin
    FpuF2iPlugin_logic_onResult_overflow = (((($signed(_zz_FpuF2iPlugin_logic_onResult_overflow) < $signed(_zz_FpuF2iPlugin_logic_onResult_overflow_2)) || (execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF)) && (! execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign)) || (execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN));
    if(when_FpuF2iPlugin_l123) begin
      FpuF2iPlugin_logic_onResult_overflow = 1'b1;
    end
  end

  assign FpuF2iPlugin_logic_onResult_underflow = ((((($signed(_zz_FpuF2iPlugin_logic_onResult_underflow) < $signed(_zz_FpuF2iPlugin_logic_onResult_underflow_2)) || ((FpuF2iPlugin_logic_onResult_signed && ($signed(_zz_FpuF2iPlugin_logic_onResult_underflow_3) == $signed(_zz_FpuF2iPlugin_logic_onResult_underflow_4))) && ((FpuF2iPlugin_logic_onResult_unsigned != FpuF2iPlugin_logic_onResult_unsignedMin) || execute_ctrl4_down_FpuF2iPlugin_logic_onShift_increment_lane0))) || ((! FpuF2iPlugin_logic_onResult_signed) && ((FpuF2iPlugin_logic_onResult_unsigned != 32'h0) || execute_ctrl4_down_FpuF2iPlugin_logic_onShift_increment_lane0))) || (execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF)) && execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign);
  assign FpuF2iPlugin_logic_onResult_isZero = (execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO);
  assign when_FpuF2iPlugin_l123 = (((((! FpuF2iPlugin_logic_onResult_i64) && (! execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign)) && execute_ctrl4_down_FpuF2iPlugin_logic_onShift_increment_lane0) && (&FpuF2iPlugin_logic_onResult_unsigned[30 : 0])) && (FpuF2iPlugin_logic_onResult_signed || FpuF2iPlugin_logic_onResult_unsigned[31]));
  always @(*) begin
    execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NV_lane0 = ((execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_quiet));
    if(!FpuF2iPlugin_logic_onResult_isZero) begin
      if(when_FpuF2iPlugin_l129) begin
        if(when_FpuF2iPlugin_l136) begin
          execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NV_lane0 = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NX_lane0 = 1'b0;
    if(!FpuF2iPlugin_logic_onResult_isZero) begin
      if(!when_FpuF2iPlugin_l129) begin
        if(when_FpuF2iPlugin_l138) begin
          execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NX_lane0 = 1'b1;
        end
      end
    end
  end

  assign when_FpuF2iPlugin_l136 = (! FpuF2iPlugin_logic_onResult_isZero);
  assign when_FpuF2iPlugin_l138 = (FpuF2iPlugin_logic_onResult_round != 2'b00);
  assign when_FpuF2iPlugin_l129 = (FpuF2iPlugin_logic_onResult_underflow || FpuF2iPlugin_logic_onResult_overflow);
  assign execute_ctrl4_down_FpuF2iPlugin_logic_onResult_RESULT_lane0 = FpuF2iPlugin_logic_onResult_resultRaw;
  assign FpuF2iPlugin_logic_iwb_valid = execute_ctrl4_down_FpuF2iPlugin_SEL_lane0;
  assign FpuF2iPlugin_logic_iwb_payload = execute_ctrl4_down_FpuF2iPlugin_logic_onResult_RESULT_lane0;
  assign FpuF2iPlugin_logic_ffwb_ats[0] = execute_ctrl4_down_FpuF2iPlugin_SEL_lane0;
  assign FpuF2iPlugin_logic_ffwb_flags_NX = execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NX_lane0;
  assign FpuF2iPlugin_logic_ffwb_flags_UF = 1'b0;
  assign FpuF2iPlugin_logic_ffwb_flags_OF = 1'b0;
  assign FpuF2iPlugin_logic_ffwb_flags_DZ = 1'b0;
  assign FpuF2iPlugin_logic_ffwb_flags_NV = execute_ctrl4_down_FpuF2iPlugin_logic_onResult_NV_lane0;
  assign FpuAddPlugin_logic_addPort_cmd_at[0] = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuAddPlugin_SEL_lane0);
  assign FpuAddPlugin_logic_addPort_cmd_rs1_mode = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode;
  assign FpuAddPlugin_logic_addPort_cmd_rs1_quiet = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet;
  assign FpuAddPlugin_logic_addPort_cmd_rs1_sign = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign;
  assign FpuAddPlugin_logic_addPort_cmd_rs1_exponent = _zz_FpuAddPlugin_logic_addPort_cmd_rs1_exponent;
  assign FpuAddPlugin_logic_addPort_cmd_rs1_mantissa = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa;
  assign FpuAddPlugin_logic_addPort_cmd_rs2_mode = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode;
  assign FpuAddPlugin_logic_addPort_cmd_rs2_quiet = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet;
  assign FpuAddPlugin_logic_addPort_cmd_rs2_exponent = _zz_FpuAddPlugin_logic_addPort_cmd_rs2_exponent;
  assign FpuAddPlugin_logic_addPort_cmd_rs2_mantissa = execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa;
  assign FpuAddPlugin_logic_addPort_cmd_rs2_sign = (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign ^ execute_ctrl2_down_FpuAddPlugin_SUB_lane0);
  assign FpuAddPlugin_logic_addPort_cmd_format = execute_ctrl2_down_FpuUtils_FORMAT_lane0;
  assign FpuAddPlugin_logic_addPort_cmd_roundMode = execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  assign FpuAddPlugin_logic_addPort_cmd_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX = 5'h0;
  assign FpuAddPlugin_logic_addPort_cmd_flags_NX = _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX[0];
  assign FpuAddPlugin_logic_addPort_cmd_flags_UF = _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX[1];
  assign FpuAddPlugin_logic_addPort_cmd_flags_OF = _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX[2];
  assign FpuAddPlugin_logic_addPort_cmd_flags_DZ = _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX[3];
  assign FpuAddPlugin_logic_addPort_cmd_flags_NV = _zz_FpuAddPlugin_logic_addPort_cmd_flags_NX[4];
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = _zz_execute_ctrl2_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_SIGN_lane0 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign ^ execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign);
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO));
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF));
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF)) && ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO)));
  assign execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN)) || execute_ctrl2_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0);
  assign FpuMulPlugin_logic_mulCmd_m1 = {1'b1,execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa};
  assign FpuMulPlugin_logic_mulCmd_m2 = {1'b1,execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa};
  assign execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0 = _zz_execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0[105 : 0];
  assign FpuMulPlugin_logic_norm_needShift = execute_ctrl5_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0[105];
  assign execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0 = _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_EXP_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0 = (FpuMulPlugin_logic_norm_needShift ? execute_ctrl5_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0[104 : 0] : _zz_execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0);
  always @(*) begin
    FpuMulPlugin_logic_onPack_nv = 1'b0;
    if(execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0) begin
      if(when_FpuMulPlugin_l148) begin
        FpuMulPlugin_logic_onPack_nv = 1'b1;
      end
    end
  end

  always @(*) begin
    FpuMulPlugin_logic_onPack_mode = FloatMode_NORMAL;
    if(execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0) begin
      FpuMulPlugin_logic_onPack_mode = FloatMode_NAN;
    end else begin
      if(execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0) begin
        FpuMulPlugin_logic_onPack_mode = FloatMode_INF;
      end else begin
        if(execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0) begin
          FpuMulPlugin_logic_onPack_mode = FloatMode_ZERO;
        end
      end
    end
  end

  assign when_FpuMulPlugin_l148 = ((execute_ctrl5_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 || ((execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_quiet))) || ((execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_quiet)));
  assign FpuMulPlugin_logic_packPort_cmd_at[0] = ((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_down_FpuMulPlugin_SEL_lane0) && (! execute_ctrl5_down_FpuMulPlugin_FMA_lane0));
  assign FpuMulPlugin_logic_packPort_cmd_value_sign = execute_ctrl5_down_FpuMulPlugin_logic_calc_SIGN_lane0;
  assign FpuMulPlugin_logic_packPort_cmd_value_exponent = _zz_FpuMulPlugin_logic_packPort_cmd_value_exponent;
  assign _zz_when_AFix_l852_1 = execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0;
  always @(*) begin
    _zz_FpuMulPlugin_logic_packPort_cmd_value_mantissa = _zz_when_AFix_l852_1[104 : 51];
    if(when_AFix_l852_1) begin
      _zz_FpuMulPlugin_logic_packPort_cmd_value_mantissa[0] = 1'b1;
    end
  end

  assign when_AFix_l852_1 = (|_zz_when_AFix_l852_1[50 : 0]);
  assign FpuMulPlugin_logic_packPort_cmd_value_mantissa = _zz_FpuMulPlugin_logic_packPort_cmd_value_mantissa;
  assign FpuMulPlugin_logic_packPort_cmd_value_mode = FpuMulPlugin_logic_onPack_mode;
  assign FpuMulPlugin_logic_packPort_cmd_value_quiet = 1'b1;
  assign FpuMulPlugin_logic_packPort_cmd_format = execute_ctrl5_down_FpuUtils_FORMAT_lane0;
  assign FpuMulPlugin_logic_packPort_cmd_roundMode = execute_ctrl5_down_FpuUtils_ROUNDING_lane0;
  assign FpuMulPlugin_logic_packPort_cmd_uopId = execute_ctrl5_down_Decode_UOP_ID_lane0;
  assign FpuMulPlugin_logic_packPort_cmd_flags_NX = 1'b0;
  assign FpuMulPlugin_logic_packPort_cmd_flags_UF = 1'b0;
  assign FpuMulPlugin_logic_packPort_cmd_flags_OF = 1'b0;
  assign FpuMulPlugin_logic_packPort_cmd_flags_DZ = 1'b0;
  assign FpuMulPlugin_logic_packPort_cmd_flags_NV = FpuMulPlugin_logic_onPack_nv;
  assign FpuMulPlugin_logic_addPort_cmd_at[0] = ((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_down_FpuMulPlugin_SEL_lane0) && execute_ctrl5_down_FpuMulPlugin_FMA_lane0);
  assign FpuMulPlugin_logic_addPort_cmd_rs1_sign = (execute_ctrl5_down_FpuMulPlugin_logic_calc_SIGN_lane0 ^ execute_ctrl5_down_FpuMulPlugin_SUB1_lane0);
  assign FpuMulPlugin_logic_addPort_cmd_rs1_exponent = _zz_FpuMulPlugin_logic_addPort_cmd_rs1_exponent;
  assign FpuMulPlugin_logic_addPort_cmd_rs1_mantissa = execute_ctrl5_down_FpuMulPlugin_logic_norm_MAN_lane0;
  assign FpuMulPlugin_logic_addPort_cmd_rs1_mode = FpuMulPlugin_logic_onPack_mode;
  assign FpuMulPlugin_logic_addPort_cmd_rs1_quiet = 1'b1;
  assign FpuMulPlugin_logic_addPort_cmd_rs2_mode = execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode;
  assign FpuMulPlugin_logic_addPort_cmd_rs2_quiet = execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_quiet;
  assign FpuMulPlugin_logic_addPort_cmd_rs2_exponent = _zz_FpuMulPlugin_logic_addPort_cmd_rs2_exponent;
  assign FpuMulPlugin_logic_addPort_cmd_rs2_mantissa = execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mantissa;
  assign FpuMulPlugin_logic_addPort_cmd_rs2_sign = (execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_sign ^ execute_ctrl5_down_FpuMulPlugin_SUB2_lane0);
  assign FpuMulPlugin_logic_addPort_cmd_format = execute_ctrl5_down_FpuUtils_FORMAT_lane0;
  assign FpuMulPlugin_logic_addPort_cmd_roundMode = execute_ctrl5_down_FpuUtils_ROUNDING_lane0;
  assign FpuMulPlugin_logic_addPort_cmd_uopId = execute_ctrl5_down_Decode_UOP_ID_lane0;
  assign FpuMulPlugin_logic_addPort_cmd_flags_NX = 1'b0;
  assign FpuMulPlugin_logic_addPort_cmd_flags_UF = 1'b0;
  assign FpuMulPlugin_logic_addPort_cmd_flags_OF = 1'b0;
  assign FpuMulPlugin_logic_addPort_cmd_flags_DZ = 1'b0;
  assign FpuMulPlugin_logic_addPort_cmd_flags_NV = FpuMulPlugin_logic_onPack_nv;
  assign when_FpuSqrtPlugin_l66 = (FpuUnpackerPlugin_logic_unpackDone && (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO));
  assign io_input_fire = (FpuSqrtPlugin_logic_sqrt_io_input_valid && FpuSqrtPlugin_logic_sqrt_io_input_ready);
  assign FpuSqrtPlugin_logic_sqrt_io_input_valid = ((((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuSqrtPlugin_SEL_lane0) && FpuUnpackerPlugin_logic_unpackDone) && (! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO))) && (! FpuSqrtPlugin_logic_onExecute_cmdSent));
  assign FpuSqrtPlugin_logic_sqrt_io_input_payload_a = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent[0] ? {{1'b1,execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa},1'b0} : {2'b01,execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa});
  assign FpuSqrtPlugin_logic_onExecute_freeze = ((((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuSqrtPlugin_SEL_lane0) && (! FpuSqrtPlugin_logic_sqrt_io_output_valid)) && (! FpuSqrtPlugin_logic_onExecute_unscheduleRequest)) && (! FpuSqrtPlugin_logic_onExecute_isZero));
  assign FpuSqrtPlugin_logic_onExecute_exp = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_exponent[11 : 1];
  assign FpuSqrtPlugin_logic_onExecute_scrap = (FpuSqrtPlugin_logic_sqrt_io_output_payload_remain != 57'h0);
  assign FpuSqrtPlugin_logic_packPort_cmd_at[0] = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuSqrtPlugin_SEL_lane0);
  assign FpuSqrtPlugin_logic_packPort_cmd_format = execute_ctrl2_down_FpuUtils_FORMAT_lane0;
  assign FpuSqrtPlugin_logic_packPort_cmd_roundMode = execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  assign FpuSqrtPlugin_logic_packPort_cmd_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  always @(*) begin
    FpuSqrtPlugin_logic_packPort_cmd_value_mode = FloatMode_NORMAL;
    if(when_FpuSqrtPlugin_l92) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_mode = FloatMode_INF;
    end
    if(FpuSqrtPlugin_logic_onExecute_negative) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_mode = FloatMode_NAN;
    end
    if(when_FpuSqrtPlugin_l101) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_mode = FloatMode_NAN;
    end
    if(when_FpuSqrtPlugin_l105) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_mode = FloatMode_ZERO;
    end
  end

  always @(*) begin
    FpuSqrtPlugin_logic_packPort_cmd_value_quiet = 1'b0;
    if(FpuSqrtPlugin_logic_onExecute_negative) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_quiet = 1'b1;
    end
    if(when_FpuSqrtPlugin_l101) begin
      FpuSqrtPlugin_logic_packPort_cmd_value_quiet = 1'b1;
    end
  end

  assign FpuSqrtPlugin_logic_packPort_cmd_value_sign = execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign;
  assign FpuSqrtPlugin_logic_packPort_cmd_value_exponent = _zz_FpuSqrtPlugin_logic_packPort_cmd_value_exponent;
  assign FpuSqrtPlugin_logic_packPort_cmd_value_mantissa = {FpuSqrtPlugin_logic_sqrt_io_output_payload_result,FpuSqrtPlugin_logic_onExecute_scrap};
  assign FpuSqrtPlugin_logic_onExecute_negative = (((! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN)) && (! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO))) && execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign);
  assign when_FpuSqrtPlugin_l92 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF);
  always @(*) begin
    FpuSqrtPlugin_logic_onExecute_NV = 1'b0;
    if(FpuSqrtPlugin_logic_onExecute_negative) begin
      FpuSqrtPlugin_logic_onExecute_NV = 1'b1;
    end
    if(when_FpuSqrtPlugin_l101) begin
      FpuSqrtPlugin_logic_onExecute_NV = (! execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet);
    end
  end

  assign when_FpuSqrtPlugin_l101 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN);
  assign when_FpuSqrtPlugin_l105 = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO);
  assign FpuSqrtPlugin_logic_packPort_cmd_flags_NX = 1'b0;
  assign FpuSqrtPlugin_logic_packPort_cmd_flags_UF = 1'b0;
  assign FpuSqrtPlugin_logic_packPort_cmd_flags_OF = 1'b0;
  assign FpuSqrtPlugin_logic_packPort_cmd_flags_DZ = 1'b0;
  assign FpuSqrtPlugin_logic_packPort_cmd_flags_NV = FpuSqrtPlugin_logic_onExecute_NV;
  assign FpuXxPlugin_logic_packPort_cmd_at[0] = (execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_down_FpuXxPlugin_SEL_lane0);
  assign _zz_FpuXxPlugin_logic_packPort_cmd_format = ((execute_ctrl3_down_FpuUtils_FORMAT_lane0 == FpuFormat_FpuCmpPlugin_logic_f32_1) ? FpuFormat_FpuCmpPlugin_logic_f64_1 : FpuFormat_FpuCmpPlugin_logic_f32_1);
  assign FpuXxPlugin_logic_packPort_cmd_format = _zz_FpuXxPlugin_logic_packPort_cmd_format;
  assign FpuXxPlugin_logic_packPort_cmd_roundMode = execute_ctrl3_down_FpuUtils_ROUNDING_lane0;
  assign FpuXxPlugin_logic_packPort_cmd_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign FpuXxPlugin_logic_packPort_cmd_value_mode = execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode;
  assign FpuXxPlugin_logic_packPort_cmd_value_sign = execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign;
  assign FpuXxPlugin_logic_packPort_cmd_value_exponent = _zz_FpuXxPlugin_logic_packPort_cmd_value_exponent;
  assign FpuXxPlugin_logic_packPort_cmd_value_mantissa = ({2'd0,execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mantissa} <<< 2'd2);
  assign FpuXxPlugin_logic_packPort_cmd_value_quiet = 1'b1;
  assign FpuXxPlugin_logic_packPort_cmd_flags_NX = 1'b0;
  assign FpuXxPlugin_logic_packPort_cmd_flags_UF = 1'b0;
  assign FpuXxPlugin_logic_packPort_cmd_flags_OF = 1'b0;
  assign FpuXxPlugin_logic_packPort_cmd_flags_DZ = 1'b0;
  assign FpuXxPlugin_logic_packPort_cmd_flags_NV = ((execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet));
  assign when_FpuDivPlugin_l68 = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuDivPlugin_SEL_lane0) && FpuUnpackerPlugin_logic_unpackDone) && (! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO)));
  assign execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0 = (early0_DivPlugin_logic_processing_div_io_rsp_payload_result[56 : 1] | _zz_execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0);
  assign FpuDivPlugin_logic_onExecute_needShift = (! execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0[55]);
  assign FpuDivPlugin_logic_onExecute_mantissa = (FpuDivPlugin_logic_onExecute_needShift ? execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0[53 : 0] : (execute_ctrl2_down_FpuDivPlugin_logic_onExecute_DIVIDER_RSP_lane0[54 : 1] | _zz_FpuDivPlugin_logic_onExecute_mantissa));
  assign FpuDivPlugin_logic_onExecute_exponent = _zz_FpuDivPlugin_logic_onExecute_exponent_1;
  assign FpuDivPlugin_logic_packPort_cmd_at[0] = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_FpuDivPlugin_SEL_lane0);
  always @(*) begin
    FpuDivPlugin_logic_packPort_cmd_value_mode = FloatMode_NORMAL;
    if(FpuDivPlugin_logic_onExecute_forceNan) begin
      FpuDivPlugin_logic_packPort_cmd_value_mode = FloatMode_NAN;
    end else begin
      if(FpuDivPlugin_logic_onExecute_forceOverflow) begin
        FpuDivPlugin_logic_packPort_cmd_value_mode = FloatMode_INF;
      end else begin
        if(FpuDivPlugin_logic_onExecute_forceZero) begin
          FpuDivPlugin_logic_packPort_cmd_value_mode = FloatMode_ZERO;
        end
      end
    end
  end

  always @(*) begin
    FpuDivPlugin_logic_packPort_cmd_value_quiet = 1'b0;
    if(FpuDivPlugin_logic_onExecute_forceNan) begin
      FpuDivPlugin_logic_packPort_cmd_value_quiet = 1'b1;
    end
  end

  assign FpuDivPlugin_logic_packPort_cmd_value_sign = (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign ^ execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign);
  assign FpuDivPlugin_logic_packPort_cmd_value_exponent = _zz_FpuDivPlugin_logic_packPort_cmd_value_exponent;
  assign FpuDivPlugin_logic_packPort_cmd_value_mantissa = FpuDivPlugin_logic_onExecute_mantissa;
  assign FpuDivPlugin_logic_packPort_cmd_format = execute_ctrl2_down_FpuUtils_FORMAT_lane0;
  assign FpuDivPlugin_logic_packPort_cmd_roundMode = execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
  assign FpuDivPlugin_logic_packPort_cmd_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign FpuDivPlugin_logic_onExecute_forceOverflow = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO));
  assign FpuDivPlugin_logic_onExecute_infinitynan = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO) && (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO)) || ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF) && (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF)));
  assign FpuDivPlugin_logic_onExecute_forceNan = (((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN)) || FpuDivPlugin_logic_onExecute_infinitynan);
  assign FpuDivPlugin_logic_onExecute_forceZero = ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_ZERO) || (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_INF));
  assign FpuDivPlugin_logic_packPort_cmd_flags_NX = 1'b0;
  assign FpuDivPlugin_logic_packPort_cmd_flags_UF = 1'b0;
  assign FpuDivPlugin_logic_packPort_cmd_flags_OF = 1'b0;
  assign FpuDivPlugin_logic_packPort_cmd_flags_DZ = (((! FpuDivPlugin_logic_onExecute_forceNan) && (! (execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_INF))) && (execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_ZERO));
  always @(*) begin
    FpuDivPlugin_logic_packPort_cmd_flags_NV = 1'b0;
    if(FpuDivPlugin_logic_onExecute_forceNan) begin
      if(when_FpuDivPlugin_l102) begin
        FpuDivPlugin_logic_packPort_cmd_flags_NV = 1'b1;
      end
    end
  end

  assign when_FpuDivPlugin_l102 = ((FpuDivPlugin_logic_onExecute_infinitynan || ((execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet))) || ((execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode == FloatMode_NAN) && (! execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet)));
  assign when_CtrlLaneApi_l50_4 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_0_fire = (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_0_decodeId = decode_ctrls_1_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOpId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOp = decode_ctrls_1_down_Decode_UOP_0;
  assign when_CtrlLaneApi_l50_5 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane1_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_1_fire = (decode_ctrls_1_up_LANE_SEL_1 && (! decode_ctrls_1_up_LANE_SEL_1_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_1_decodeId = decode_ctrls_1_down_Decode_DOP_ID_1;
  assign WhiteboxerPlugin_logic_serializeds_1_microOpId = decode_ctrls_1_down_Decode_UOP_ID_1;
  assign WhiteboxerPlugin_logic_serializeds_1_microOp = decode_ctrls_1_down_Decode_UOP_1;
  assign when_CtrlLaneApi_l50_6 = (execute_ctrl0_down_isReady || execute_lane0_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_0_fire = (execute_ctrl0_down_LANE_SEL_lane0 && (! execute_ctrl0_down_LANE_SEL_lane0_regNext));
  assign WhiteboxerPlugin_logic_dispatches_0_microOpId = execute_ctrl0_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l50_7 = (execute_ctrl0_down_isReady || execute_lane1_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_1_fire = (execute_ctrl0_down_LANE_SEL_lane1 && (! execute_ctrl0_down_LANE_SEL_lane1_regNext));
  assign WhiteboxerPlugin_logic_dispatches_1_microOpId = execute_ctrl0_down_Decode_UOP_ID_lane1;
  assign when_CtrlLaneApi_l50_8 = (execute_ctrl2_down_isReady || execute_lane0_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_0_fire = ((execute_ctrl2_down_LANE_SEL_lane0 && (! execute_ctrl2_down_LANE_SEL_lane0_regNext)) && execute_ctrl2_down_COMMIT_lane0);
  assign WhiteboxerPlugin_logic_executes_0_microOpId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l50_9 = (execute_ctrl2_down_isReady || execute_lane1_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_1_fire = ((execute_ctrl2_down_LANE_SEL_lane1 && (! execute_ctrl2_down_LANE_SEL_lane1_regNext)) && execute_ctrl2_down_COMMIT_lane1);
  assign WhiteboxerPlugin_logic_executes_1_microOpId = execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign BtbPlugin_logic_onForget_hash = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[21 : 10];
  assign BtbPlugin_logic_memRead_cmd_valid = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_memRead_cmd_payload = _zz_BtbPlugin_logic_memRead_cmd_payload[6:0];
  assign fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS = ((BtbPlugin_logic_memWrite_valid && (BtbPlugin_logic_memWrite_payload_address == BtbPlugin_logic_memRead_cmd_payload)) ? BtbPlugin_logic_memWrite_payload_mask : 2'b00);
  assign fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200 = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_predictions = {fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3[1],{fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2[1],{fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1[1],fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[1]}}};
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash = BtbPlugin_logic_memRead_rsp_0_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow = BtbPlugin_logic_memRead_rsp_0_sliceLow;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget = BtbPlugin_logic_memRead_rsp_0_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch = BtbPlugin_logic_memRead_rsp_0_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush = BtbPlugin_logic_memRead_rsp_0_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop = BtbPlugin_logic_memRead_rsp_0_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 10]) && (fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 1] <= {1'b0,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow}));
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN = ((! fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[{1'b0,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow}]);
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash = BtbPlugin_logic_memRead_rsp_1_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow = BtbPlugin_logic_memRead_rsp_1_sliceLow;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget = BtbPlugin_logic_memRead_rsp_1_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch = BtbPlugin_logic_memRead_rsp_1_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush = BtbPlugin_logic_memRead_rsp_1_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop = BtbPlugin_logic_memRead_rsp_1_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 10]) && (fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 1] <= {1'b1,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow}));
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN = ((! fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[{1'b1,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow}]);
  assign BtbPlugin_logic_ras_readIt = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_applyIt_chunksMask = {(fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN) == 1'b0)),(fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && 1'b1)};
  assign BtbPlugin_logic_applyIt_chunksTakenOh = ({fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN} & BtbPlugin_logic_applyIt_chunksMask);
  assign BtbPlugin_logic_applyIt_needIt = (fetch_logic_ctrls_1_up_isValid && (|BtbPlugin_logic_applyIt_chunksTakenOh));
  assign when_BtbPlugin_l233 = (fetch_logic_ctrls_1_up_isReady || fetch_logic_ctrls_1_up_isCancel);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign _zz_BtbPlugin_logic_applyIt_doItSlice = BtbPlugin_logic_applyIt_chunksTakenOh[1];
  assign _zz_BtbPlugin_logic_applyIt_entry_hash = ((BtbPlugin_logic_applyIt_chunksTakenOh[0] ? {fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop,{fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush,{fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch,{_zz__zz_BtbPlugin_logic_applyIt_entry_hash,_zz__zz_BtbPlugin_logic_applyIt_entry_hash_1}}}} : 47'h0) | (_zz_BtbPlugin_logic_applyIt_doItSlice ? {fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop,{fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush,{fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch,{_zz__zz_BtbPlugin_logic_applyIt_entry_hash_2,_zz__zz_BtbPlugin_logic_applyIt_entry_hash_3}}}} : 47'h0));
  assign BtbPlugin_logic_applyIt_entry_hash = _zz_BtbPlugin_logic_applyIt_entry_hash[11 : 0];
  assign BtbPlugin_logic_applyIt_entry_sliceLow = _zz_BtbPlugin_logic_applyIt_entry_hash[12 : 12];
  assign BtbPlugin_logic_applyIt_entry_pcTarget = _zz_BtbPlugin_logic_applyIt_entry_hash[43 : 13];
  assign BtbPlugin_logic_applyIt_entry_isBranch = _zz_BtbPlugin_logic_applyIt_entry_hash[44];
  assign BtbPlugin_logic_applyIt_entry_isPush = _zz_BtbPlugin_logic_applyIt_entry_hash[45];
  assign BtbPlugin_logic_applyIt_entry_isPop = _zz_BtbPlugin_logic_applyIt_entry_hash[46];
  always @(*) begin
    BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_applyIt_entry_pcTarget;
    if(BtbPlugin_logic_applyIt_entry_isPop) begin
      BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_ras_read;
    end
  end

  assign BtbPlugin_logic_applyIt_doItSlice = {_zz_BtbPlugin_logic_applyIt_doItSlice,BtbPlugin_logic_applyIt_entry_sliceLow};
  assign BtbPlugin_logic_applyIt_rasLogic_pushValid = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPush);
  always @(*) begin
    BtbPlugin_logic_applyIt_rasLogic_pushPc = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
    BtbPlugin_logic_applyIt_rasLogic_pushPc[2 : 1] = BtbPlugin_logic_applyIt_doItSlice;
  end

  assign when_BtbPlugin_l246 = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPop);
  assign BtbPlugin_logic_flushPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_flushPort_payload_self = 1'b0;
  assign BtbPlugin_logic_pcPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_pcPort_payload_fault = 1'b0;
  assign BtbPlugin_logic_pcPort_payload_pc = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED = BtbPlugin_logic_applyIt_needIt;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE = BtbPlugin_logic_applyIt_doItSlice;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign BtbPlugin_logic_applyIt_history_layers_0_history = fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_doIt = (BtbPlugin_logic_applyIt_chunksMask[0] && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_shifted = {BtbPlugin_logic_applyIt_history_layers_0_history[10 : 0],fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_1_history = (BtbPlugin_logic_applyIt_history_layersLogic_0_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_0_shifted : BtbPlugin_logic_applyIt_history_layers_0_history);
  assign BtbPlugin_logic_applyIt_history_layersLogic_1_doIt = (BtbPlugin_logic_applyIt_chunksMask[1] && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_1_shifted = {BtbPlugin_logic_applyIt_history_layers_1_history[10 : 0],fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_2_history = (BtbPlugin_logic_applyIt_history_layersLogic_1_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_1_shifted : BtbPlugin_logic_applyIt_history_layers_1_history);
  assign BtbPlugin_logic_historyPort_valid = ((fetch_logic_ctrls_1_up_isValid && (! BtbPlugin_logic_applyIt_correctionSent)) && (|{fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT}));
  assign BtbPlugin_logic_historyPort_payload_history = BtbPlugin_logic_applyIt_history_layers_2_history;
  always @(*) begin
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[0] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b0));
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[1] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b1));
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[2] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow == 1'b0));
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[3] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow == 1'b1));
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[0] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[1] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[2] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[3] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
  end

  assign AlignerPlugin_logic_buffer_flushIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && _zz_AlignerPlugin_logic_buffer_flushIt),{_zz_AlignerPlugin_logic_buffer_flushIt_1,{_zz_AlignerPlugin_logic_buffer_flushIt_2,_zz_AlignerPlugin_logic_buffer_flushIt_3}}}}}}});
  assign AlignerPlugin_logic_buffer_readers_0_firstFromBuffer = (|{_zz_AlignerPlugin_logic_extractors_0_redo_3,{_zz_AlignerPlugin_logic_extractors_0_redo_2,{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo}}});
  assign AlignerPlugin_logic_buffer_readers_0_lastFromBuffer = ({AlignerPlugin_logic_extractors_0_usageMask[7],{AlignerPlugin_logic_extractors_0_usageMask[6],{AlignerPlugin_logic_extractors_0_usageMask[5],AlignerPlugin_logic_extractors_0_usageMask[4]}}} == 4'b0000);
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction = {_zz_AlignerPlugin_logic_extractors_0_redo_7,{_zz_AlignerPlugin_logic_extractors_0_redo_6,{_zz_AlignerPlugin_logic_extractors_0_redo_5,{_zz_AlignerPlugin_logic_extractors_0_redo_4,{_zz_AlignerPlugin_logic_extractors_0_redo_3,{_zz_AlignerPlugin_logic_extractors_0_redo_2,{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo}}}}}}};
  assign AlignerPlugin_logic_extractors_0_ctx_instruction = ((((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1 ? AlignerPlugin_logic_slicesInstructions_0 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3 ? AlignerPlugin_logic_slicesInstructions_1 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4)) | ((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5 ? AlignerPlugin_logic_slicesInstructions_2 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7 ? AlignerPlugin_logic_slicesInstructions_3 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8))) | (((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9 ? AlignerPlugin_logic_slicesInstructions_4 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11 ? AlignerPlugin_logic_slicesInstructions_5 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12)) | ((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13 ? AlignerPlugin_logic_slicesInstructions_6 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15 ? AlignerPlugin_logic_slicesInstructions_7 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16))));
  always @(*) begin
    AlignerPlugin_logic_extractors_0_ctx_pc = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_pc : fetch_logic_ctrls_2_down_Fetch_WORD_PC);
    AlignerPlugin_logic_extractors_0_ctx_pc[2 : 1] = {_zz_AlignerPlugin_logic_extractors_0_ctx_pc_2,_zz_AlignerPlugin_logic_extractors_0_ctx_pc_1};
  end

  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc = (|{_zz_AlignerPlugin_logic_extractors_0_redo_7,_zz_AlignerPlugin_logic_extractors_0_redo_3});
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc_1 = ((|{_zz_AlignerPlugin_logic_extractors_0_redo_5,_zz_AlignerPlugin_logic_extractors_0_redo_1}) || _zz_AlignerPlugin_logic_extractors_0_ctx_pc);
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc_2 = ((|{_zz_AlignerPlugin_logic_extractors_0_redo_6,_zz_AlignerPlugin_logic_extractors_0_redo_2}) || _zz_AlignerPlugin_logic_extractors_0_ctx_pc);
  assign AlignerPlugin_logic_extractors_0_ctx_trap = ((AlignerPlugin_logic_buffer_readers_0_firstFromBuffer && AlignerPlugin_logic_buffer_trap) || ((! AlignerPlugin_logic_buffer_readers_0_lastFromBuffer) && fetch_logic_ctrls_2_down_TRAP));
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_hm_Fetch_ID : fetch_logic_ctrls_2_down_Fetch_ID);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY : fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED : fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign AlignerPlugin_logic_buffer_readers_1_firstFromBuffer = (|{_zz_AlignerPlugin_logic_extractors_1_redo_2,{_zz_AlignerPlugin_logic_extractors_1_redo_1,_zz_AlignerPlugin_logic_extractors_1_redo}});
  assign AlignerPlugin_logic_buffer_readers_1_lastFromBuffer = ({AlignerPlugin_logic_extractors_1_usageMask[7],{AlignerPlugin_logic_extractors_1_usageMask[6],{AlignerPlugin_logic_extractors_1_usageMask[5],AlignerPlugin_logic_extractors_1_usageMask[4]}}} == 4'b0000);
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_instruction = {_zz_AlignerPlugin_logic_extractors_1_redo_6,{_zz_AlignerPlugin_logic_extractors_1_redo_5,{_zz_AlignerPlugin_logic_extractors_1_redo_4,{_zz_AlignerPlugin_logic_extractors_1_redo_3,{_zz_AlignerPlugin_logic_extractors_1_redo_2,{_zz_AlignerPlugin_logic_extractors_1_redo_1,_zz_AlignerPlugin_logic_extractors_1_redo}}}}}};
  assign AlignerPlugin_logic_extractors_1_ctx_instruction = ((((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[0] ? AlignerPlugin_logic_slicesInstructions_1 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[1] ? AlignerPlugin_logic_slicesInstructions_2 : 32'h0)) | ((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[2] ? AlignerPlugin_logic_slicesInstructions_3 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[3] ? AlignerPlugin_logic_slicesInstructions_4 : 32'h0))) | (((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[4] ? AlignerPlugin_logic_slicesInstructions_5 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[5] ? AlignerPlugin_logic_slicesInstructions_6 : 32'h0)) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[6] ? AlignerPlugin_logic_slicesInstructions_7 : 32'h0)));
  always @(*) begin
    AlignerPlugin_logic_extractors_1_ctx_pc = (AlignerPlugin_logic_buffer_readers_1_firstFromBuffer ? AlignerPlugin_logic_buffer_pc : fetch_logic_ctrls_2_down_Fetch_WORD_PC);
    AlignerPlugin_logic_extractors_1_ctx_pc[2 : 1] = {_zz_AlignerPlugin_logic_extractors_1_ctx_pc_2,_zz_AlignerPlugin_logic_extractors_1_ctx_pc_1};
  end

  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc = (|{_zz_AlignerPlugin_logic_extractors_1_redo_6,_zz_AlignerPlugin_logic_extractors_1_redo_2});
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc_1 = ((|{_zz_AlignerPlugin_logic_extractors_1_redo_4,_zz_AlignerPlugin_logic_extractors_1_redo}) || _zz_AlignerPlugin_logic_extractors_1_ctx_pc);
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc_2 = ((|{_zz_AlignerPlugin_logic_extractors_1_redo_5,_zz_AlignerPlugin_logic_extractors_1_redo_1}) || _zz_AlignerPlugin_logic_extractors_1_ctx_pc);
  assign AlignerPlugin_logic_extractors_1_ctx_trap = ((AlignerPlugin_logic_buffer_readers_1_firstFromBuffer && AlignerPlugin_logic_buffer_trap) || ((! AlignerPlugin_logic_buffer_readers_1_lastFromBuffer) && fetch_logic_ctrls_2_down_TRAP));
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID = (AlignerPlugin_logic_buffer_readers_1_firstFromBuffer ? AlignerPlugin_logic_buffer_hm_Fetch_ID : fetch_logic_ctrls_2_down_Fetch_ID);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY : fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED : fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign AlignerPlugin_api_downMoving = decode_ctrls_0_up_isMoving;
  assign DispatchPlugin_logic_candidates_0_cancel = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && _zz_DispatchPlugin_logic_candidates_0_cancel),(LsuPlugin_logic_flushPort_valid && _zz_DispatchPlugin_logic_candidates_0_cancel_1)}}}}}});
  assign DispatchPlugin_logic_slotsFeeds_free = (&DispatchPlugin_logic_candidates_0_moving);
  assign DispatchPlugin_logic_slotsFeeds_fit = (_zz_DispatchPlugin_logic_slotsFeeds_fit <= 2'b01);
  assign DispatchPlugin_logic_slotsFeeds_doIt = (DispatchPlugin_logic_slotsFeeds_free && DispatchPlugin_logic_slotsFeeds_fit);
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid = {(! DispatchPlugin_logic_candidates_2_moving),(! DispatchPlugin_logic_candidates_1_moving)};
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_1 = _zz_DispatchPlugin_logic_slots_0_ctx_valid[0];
  always @(*) begin
    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2[0] = (_zz_DispatchPlugin_logic_slots_0_ctx_valid_1 && (! 1'b0));
    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2[1] = (_zz_DispatchPlugin_logic_slots_0_ctx_valid[1] && (! _zz_DispatchPlugin_logic_slots_0_ctx_valid_1));
  end

  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_3 = _zz_DispatchPlugin_logic_slots_0_ctx_valid_2;
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_4 = ((_zz_DispatchPlugin_logic_slots_0_ctx_valid_3[0] ? {{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1}},{DispatchPlugin_logic_candidates_1_ctx_uop,{DispatchPlugin_logic_candidates_1_ctx_laneLayerHits,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14}}} : 198'h0) | (_zz_DispatchPlugin_logic_slots_0_ctx_valid_3[1] ? {{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16}},{DispatchPlugin_logic_candidates_2_ctx_uop,{DispatchPlugin_logic_candidates_2_ctx_laneLayerHits,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_29}}} : 198'h0));
  assign _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED = _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[197 : 37];
  assign _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[48 : 41];
  assign DispatchPlugin_logic_scheduler_eusFree_0 = 2'b11;
  assign DispatchPlugin_logic_scheduler_hartFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_arbiters_0_candHazard = 1'b0;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits = (((DispatchPlugin_logic_candidates_0_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_0_rsHazards)) & (~ DispatchPlugin_logic_candidates_0_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_0[0],{DispatchPlugin_logic_scheduler_eusFree_0[1],{DispatchPlugin_logic_scheduler_eusFree_0[0],DispatchPlugin_logic_scheduler_eusFree_0[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_0_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_0_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_0_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_0_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_0_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_0_doIt = (((((DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_flushHazards)) && (! DispatchPlugin_logic_candidates_0_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_0[0]) && (! DispatchPlugin_logic_scheduler_arbiters_0_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_1 = (DispatchPlugin_logic_scheduler_eusFree_0 & ((! DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_0_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_1 = (DispatchPlugin_logic_scheduler_hartFree_0 & (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_0_fire = ((DispatchPlugin_logic_scheduler_arbiters_0_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite = ((DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_3 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RS3_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit = (DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_3,{DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1,DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0}}}));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazard = (|DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit);
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits = (((DispatchPlugin_logic_candidates_1_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_1_rsHazards)) & (~ DispatchPlugin_logic_candidates_1_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_1[0],{DispatchPlugin_logic_scheduler_eusFree_1[1],{DispatchPlugin_logic_scheduler_eusFree_1[0],DispatchPlugin_logic_scheduler_eusFree_1[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_1_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_1_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_1_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_1_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_1_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_1_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_1_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_1_doIt = (((((DispatchPlugin_logic_candidates_1_ctx_valid && (! DispatchPlugin_logic_candidates_1_flushHazards)) && (! DispatchPlugin_logic_candidates_1_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_1_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_1[0]) && (! DispatchPlugin_logic_scheduler_arbiters_1_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_2 = (DispatchPlugin_logic_scheduler_eusFree_1 & ((! DispatchPlugin_logic_scheduler_arbiters_1_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_1_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_2 = (DispatchPlugin_logic_scheduler_hartFree_1 & (((! DispatchPlugin_logic_candidates_1_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_1_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_1_fire = ((DispatchPlugin_logic_scheduler_arbiters_1_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite = ((DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_3 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit = (DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_3,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0}}}));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite = ((DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS)) && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_3 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS3_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS)) && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID == DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit = (DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_3,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0}}}));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazard = (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits = (((DispatchPlugin_logic_candidates_2_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_2_rsHazards)) & (~ DispatchPlugin_logic_candidates_2_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_2[0],{DispatchPlugin_logic_scheduler_eusFree_2[1],{DispatchPlugin_logic_scheduler_eusFree_2[0],DispatchPlugin_logic_scheduler_eusFree_2[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_2_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_2_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_2_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_2_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_2_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_2_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_2_doIt = (((((DispatchPlugin_logic_candidates_2_ctx_valid && (! DispatchPlugin_logic_candidates_2_flushHazards)) && (! DispatchPlugin_logic_candidates_2_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_2_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_2[0]) && (! DispatchPlugin_logic_scheduler_arbiters_2_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_3 = (DispatchPlugin_logic_scheduler_eusFree_2 & ((! DispatchPlugin_logic_scheduler_arbiters_2_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_2_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_3 = (DispatchPlugin_logic_scheduler_hartFree_2 & (((! DispatchPlugin_logic_candidates_2_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_2_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_2_fire = ((DispatchPlugin_logic_scheduler_arbiters_2_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_inserter_0_oh = {(DispatchPlugin_logic_scheduler_arbiters_2_doIt && DispatchPlugin_logic_scheduler_arbiters_2_eusOh[0]),{(DispatchPlugin_logic_scheduler_arbiters_1_doIt && DispatchPlugin_logic_scheduler_arbiters_1_eusOh[0]),(DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[0])}};
  assign _zz_execute_ctrl0_up_LANE_AGE_lane0 = DispatchPlugin_logic_inserter_0_oh[0];
  assign _zz_execute_ctrl0_up_LANE_AGE_lane0_1 = DispatchPlugin_logic_inserter_0_oh[1];
  assign _zz_execute_ctrl0_up_LANE_AGE_lane0_2 = DispatchPlugin_logic_inserter_0_oh[2];
  assign DispatchPlugin_logic_inserter_0_trap = _zz_DispatchPlugin_logic_inserter_0_trap[0];
  assign execute_ctrl0_up_LANE_SEL_lane0 = (((|DispatchPlugin_logic_inserter_0_oh) && (! _zz_execute_ctrl0_up_LANE_SEL_lane0[0])) && (! DispatchPlugin_api_haltDispatch));
  assign execute_ctrl0_up_Decode_UOP_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_uop : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_uop : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_uop : 32'h0));
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0[0];
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0));
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000));
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000));
  assign _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0,_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1}} : 8'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2,_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3}} : 8'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4,_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5}}} : 8'h0));
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[1 : 0];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[3 : 2];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[5 : 4];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[7 : 6];
  assign execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0));
  assign execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0[0];
  always @(*) begin
    execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0[0];
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0[0];
  assign execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0));
  assign execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane0 = _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane0[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0[0];
  assign execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane0 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane0[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0[0];
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0[0];
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0[0];
  assign execute_ctrl0_up_PC_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_PC : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_PC : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_PC : 32'h0));
  assign execute_ctrl0_up_TRAP_lane0 = _zz_execute_ctrl0_up_TRAP_lane0[0];
  assign execute_ctrl0_up_Decode_UOP_ID_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID : 16'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID : 16'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID : 16'h0));
  assign execute_ctrl0_up_RS1_ENABLE_lane0 = _zz_execute_ctrl0_up_RS1_ENABLE_lane0[0];
  assign execute_ctrl0_up_RS1_RFID_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID : 1'b0));
  assign execute_ctrl0_up_RS1_PHYS_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS : 5'h0));
  assign execute_ctrl0_up_RS2_ENABLE_lane0 = _zz_execute_ctrl0_up_RS2_ENABLE_lane0[0];
  assign execute_ctrl0_up_RS2_RFID_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID : 1'b0));
  assign execute_ctrl0_up_RS2_PHYS_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS : 5'h0));
  always @(*) begin
    execute_ctrl0_up_RD_ENABLE_lane0 = _zz_execute_ctrl0_up_RD_ENABLE_lane0[0];
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_RD_ENABLE_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_RD_RFID_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID : 1'b0));
  assign execute_ctrl0_up_RD_PHYS_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS : 5'h0));
  assign execute_ctrl0_up_RS3_ENABLE_lane0 = _zz_execute_ctrl0_up_RS3_ENABLE_lane0[0];
  assign execute_ctrl0_up_RS3_RFID_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID : 1'b0));
  assign execute_ctrl0_up_RS3_PHYS_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS : 5'h0));
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0[0];
  assign when_DispatchPlugin_l439 = ((! execute_ctrl0_up_LANE_SEL_lane0) || DispatchPlugin_logic_inserter_0_trap);
  assign execute_ctrl0_up_LANE_AGE_lane0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_age : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_age : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_age : 1'b0));
  assign execute_ctrl0_up_COMPLETED_lane0 = DispatchPlugin_logic_inserter_0_trap;
  assign DispatchPlugin_logic_inserter_0_layerOhUnfiltred = (((_zz_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_scheduler_arbiters_1_layerOh : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_scheduler_arbiters_2_layerOh : 4'b0000));
  assign DispatchPlugin_logic_inserter_0_layer_0_0 = 1'b1;
  assign DispatchPlugin_logic_inserter_0_layer_0_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[1];
  assign DispatchPlugin_logic_inserter_0_layer_1_0 = 1'b0;
  assign DispatchPlugin_logic_inserter_0_layer_1_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[3];
  assign _zz_execute_ctrl0_up_lane0_LAYER_SEL_lane0 = {DispatchPlugin_logic_inserter_0_layer_1_1,DispatchPlugin_logic_inserter_0_layer_0_1};
  assign execute_ctrl0_up_lane0_LAYER_SEL_lane0 = ((_zz_execute_ctrl0_up_lane0_LAYER_SEL_lane0[0] ? DispatchPlugin_logic_inserter_0_layer_0_0 : 1'b0) | (_zz_execute_ctrl0_up_lane0_LAYER_SEL_lane0[1] ? DispatchPlugin_logic_inserter_0_layer_1_0 : 1'b0));
  assign DispatchPlugin_logic_inserter_1_oh = {(DispatchPlugin_logic_scheduler_arbiters_2_doIt && DispatchPlugin_logic_scheduler_arbiters_2_eusOh[1]),{(DispatchPlugin_logic_scheduler_arbiters_1_doIt && DispatchPlugin_logic_scheduler_arbiters_1_eusOh[1]),(DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[1])}};
  assign _zz_execute_ctrl0_up_LANE_AGE_lane1 = DispatchPlugin_logic_inserter_1_oh[0];
  assign _zz_execute_ctrl0_up_LANE_AGE_lane1_1 = DispatchPlugin_logic_inserter_1_oh[1];
  assign _zz_execute_ctrl0_up_LANE_AGE_lane1_2 = DispatchPlugin_logic_inserter_1_oh[2];
  assign DispatchPlugin_logic_inserter_1_trap = _zz_DispatchPlugin_logic_inserter_1_trap[0];
  assign execute_ctrl0_up_LANE_SEL_lane1 = (((|DispatchPlugin_logic_inserter_1_oh) && (! _zz_execute_ctrl0_up_LANE_SEL_lane1[0])) && (! DispatchPlugin_api_haltDispatch));
  assign execute_ctrl0_up_Decode_UOP_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_uop : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_uop : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_uop : 32'h0));
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1 = _zz_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1[0];
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0));
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000));
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000));
  assign _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0,_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1}}} : 8'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2,_zz__zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3}}} : 8'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}} : 8'h0));
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[1 : 0];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[3 : 2];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[5 : 4];
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3 = _zz_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[7 : 6];
  assign execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0));
  assign execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1[0];
  always @(*) begin
    execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1[0];
    if(when_DispatchPlugin_l439_1) begin
      execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = 1'b0;
    end
  end

  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1[0];
  assign execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0));
  assign execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane1 = _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2_lane1[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane1 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane1[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane1 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane1[0];
  assign execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane1 = _zz_execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane1[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane1 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane1[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane1 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_2_lane1[0];
  assign execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane1 = _zz_execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane1[0];
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1 = _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1[0];
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1 = _zz_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1[0];
  assign execute_ctrl0_up_PC_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_PC : 32'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_PC : 32'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_PC : 32'h0));
  assign execute_ctrl0_up_TRAP_lane1 = _zz_execute_ctrl0_up_TRAP_lane1[0];
  assign execute_ctrl0_up_Decode_UOP_ID_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID : 16'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID : 16'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID : 16'h0));
  assign execute_ctrl0_up_RS1_ENABLE_lane1 = _zz_execute_ctrl0_up_RS1_ENABLE_lane1[0];
  assign execute_ctrl0_up_RS1_RFID_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_RFID : 1'b0));
  assign execute_ctrl0_up_RS1_PHYS_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS : 5'h0));
  assign execute_ctrl0_up_RS2_ENABLE_lane1 = _zz_execute_ctrl0_up_RS2_ENABLE_lane1[0];
  assign execute_ctrl0_up_RS2_RFID_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_RFID : 1'b0));
  assign execute_ctrl0_up_RS2_PHYS_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS : 5'h0));
  always @(*) begin
    execute_ctrl0_up_RD_ENABLE_lane1 = _zz_execute_ctrl0_up_RD_ENABLE_lane1[0];
    if(when_DispatchPlugin_l439_1) begin
      execute_ctrl0_up_RD_ENABLE_lane1 = 1'b0;
    end
  end

  assign execute_ctrl0_up_RD_RFID_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_RFID : 1'b0));
  assign execute_ctrl0_up_RD_PHYS_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS : 5'h0));
  assign execute_ctrl0_up_RS3_ENABLE_lane1 = _zz_execute_ctrl0_up_RS3_ENABLE_lane1[0];
  assign execute_ctrl0_up_RS3_RFID_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_RFID : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_RFID : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_RFID : 1'b0));
  assign execute_ctrl0_up_RS3_PHYS_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS3_PHYS : 5'h0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS3_PHYS : 5'h0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS3_PHYS : 5'h0));
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1[0];
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1 = _zz_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1[0];
  assign when_DispatchPlugin_l439_1 = ((! execute_ctrl0_up_LANE_SEL_lane1) || DispatchPlugin_logic_inserter_1_trap);
  assign execute_ctrl0_up_LANE_AGE_lane1 = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_age : 1'b0) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_age : 1'b0)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_age : 1'b0));
  assign execute_ctrl0_up_COMPLETED_lane1 = DispatchPlugin_logic_inserter_1_trap;
  assign DispatchPlugin_logic_inserter_1_layerOhUnfiltred = (((_zz_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 4'b0000) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_scheduler_arbiters_1_layerOh : 4'b0000)) | (_zz_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_scheduler_arbiters_2_layerOh : 4'b0000));
  assign DispatchPlugin_logic_inserter_1_layer_0_0 = 1'b1;
  assign DispatchPlugin_logic_inserter_1_layer_0_1 = DispatchPlugin_logic_inserter_1_layerOhUnfiltred[0];
  assign DispatchPlugin_logic_inserter_1_layer_1_0 = 1'b0;
  assign DispatchPlugin_logic_inserter_1_layer_1_1 = DispatchPlugin_logic_inserter_1_layerOhUnfiltred[2];
  assign _zz_execute_ctrl0_up_lane1_LAYER_SEL_lane1 = {DispatchPlugin_logic_inserter_1_layer_1_1,DispatchPlugin_logic_inserter_1_layer_0_1};
  assign execute_ctrl0_up_lane1_LAYER_SEL_lane1 = ((_zz_execute_ctrl0_up_lane1_LAYER_SEL_lane1[0] ? DispatchPlugin_logic_inserter_1_layer_0_0 : 1'b0) | (_zz_execute_ctrl0_up_lane1_LAYER_SEL_lane1[1] ? DispatchPlugin_logic_inserter_1_layer_1_0 : 1'b0));
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_address = 2'bxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = 2'b11;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = 2'b01;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign decode_logic_flushes_0_onLanes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_0_onLanes_0_doIt),{_zz_decode_logic_flushes_0_onLanes_0_doIt_1,{_zz_decode_logic_flushes_0_onLanes_0_doIt_2,_zz_decode_logic_flushes_0_onLanes_0_doIt_3}}}}}}}});
  assign decode_ctrls_0_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_0_lane0_upIsCancel = decode_logic_flushes_0_onLanes_0_doIt;
  assign decode_logic_flushes_0_onLanes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_0_onLanes_1_doIt),{_zz_decode_logic_flushes_0_onLanes_1_doIt_1,{_zz_decode_logic_flushes_0_onLanes_1_doIt_2,_zz_decode_logic_flushes_0_onLanes_1_doIt_3}}}}}}}});
  assign decode_ctrls_0_lane1_downIsCancel = 1'b0;
  assign decode_ctrls_0_lane1_upIsCancel = decode_logic_flushes_0_onLanes_1_doIt;
  assign decode_logic_flushes_1_onLanes_0_doIt = (|{((DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_0_doIt) || (_zz_decode_logic_flushes_1_onLanes_0_doIt_1 && DecoderPlugin_logic_laneLogic_1_flushPort_payload_self))),{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_0_doIt_2) && (_zz_decode_logic_flushes_1_onLanes_0_doIt_3 || _zz_decode_logic_flushes_1_onLanes_0_doIt_4)),{(late1_BranchPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_0_doIt_5),{_zz_decode_logic_flushes_1_onLanes_0_doIt_6,{_zz_decode_logic_flushes_1_onLanes_0_doIt_7,_zz_decode_logic_flushes_1_onLanes_0_doIt_8}}}}});
  assign decode_ctrls_1_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_1_lane0_upIsCancel = decode_logic_flushes_1_onLanes_0_doIt;
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt = 1'b1;
  assign decode_logic_flushes_1_onLanes_1_doIt = (|{((DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_1_doIt) || ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge == _zz_decode_logic_flushes_1_onLanes_1_doIt) && DecoderPlugin_logic_laneLogic_1_flushPort_payload_self))),{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_1_doIt) || (_zz_decode_logic_flushes_1_onLanes_1_doIt_1 && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self))),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_1_doIt_2),{_zz_decode_logic_flushes_1_onLanes_1_doIt_3,{_zz_decode_logic_flushes_1_onLanes_1_doIt_4,_zz_decode_logic_flushes_1_onLanes_1_doIt_5}}}}}});
  assign decode_ctrls_1_lane1_downIsCancel = 1'b0;
  assign decode_ctrls_1_lane1_upIsCancel = decode_logic_flushes_1_onLanes_1_doIt;
  assign decode_logic_trapPending[0] = (|{((decode_ctrls_1_up_LANE_SEL_1 && 1'b1) && decode_ctrls_1_down_TRAP_1),{((decode_ctrls_1_up_LANE_SEL_0 && 1'b1) && decode_ctrls_1_down_TRAP_0),{((decode_ctrls_0_up_LANE_SEL_1 && 1'b1) && decode_ctrls_0_down_TRAP_1),((decode_ctrls_0_up_LANE_SEL_0 && 1'b1) && decode_ctrls_0_down_TRAP_0)}}});
  assign execute_lane1_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign execute_lane1_bypasser_integer_RS1_port_address = execute_ctrl0_down_RS1_PHYS_lane1[4 : 0];
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_address = 2'bxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = 2'b01;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = 2'b10;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
        if(TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg) begin
          TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_valid = 1'b0;
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_code = 4'bxxxx;
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0111;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0011;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1011;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'bxx;
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
    end
  end

  assign when_TrapPlugin_l201 = (PrivilegedPlugin_logic_harts_0_m_status_mie || (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege));
  assign when_TrapPlugin_l207 = ((_zz_when_TrapPlugin_l207 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l207_1 = ((_zz_when_TrapPlugin_l207_1 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l207_2 = ((_zz_when_TrapPlugin_l207_2 && 1'b1) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_interrupt_pendingInterrupt = (TrapPlugin_logic_harts_0_interrupt_validBuffer && PrivilegedPlugin_api_harts_0_allowInterrupts);
  assign when_TrapPlugin_l226 = (|{_zz_when_TrapPlugin_l207_2,{_zz_when_TrapPlugin_l207_1,_zz_when_TrapPlugin_l207}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (early0_EnvPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (FetchL1Plugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (LsuPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 = (CsrAccessPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (DecoderPlugin_logic_laneLogic_0_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 = (DecoderPlugin_logic_laneLogic_1_trapPort_valid && 1'b1);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception = LsuPlugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval = LsuPlugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code = LsuPlugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg = LsuPlugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && (early0_EnvPlugin_logic_trapPort_payload_laneAge < CsrAccessPlugin_logic_trapPort_payload_laneAge))))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && (CsrAccessPlugin_logic_trapPort_payload_laneAge < early0_EnvPlugin_logic_trapPort_payload_laneAge)))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[0] ? {early0_EnvPlugin_logic_trapPort_payload_arg,{early0_EnvPlugin_logic_trapPort_payload_code,{early0_EnvPlugin_logic_trapPort_payload_tval,early0_EnvPlugin_logic_trapPort_payload_exception}}} : 39'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[1] ? {CsrAccessPlugin_logic_trapPort_payload_arg,{CsrAccessPlugin_logic_trapPort_payload_code,{CsrAccessPlugin_logic_trapPort_payload_tval,CsrAccessPlugin_logic_trapPort_payload_exception}}} : 39'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[38 : 37];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && (DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge < DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge))))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && (DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge < DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge)))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[0] ? {DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg,{DecoderPlugin_logic_laneLogic_0_trapPort_payload_code,{DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval,DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception}}} : 39'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[1] ? {DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg,{DecoderPlugin_logic_laneLogic_1_trapPort_payload_code,{DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval,DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception}}} : 39'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[38 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception = FetchL1Plugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval = FetchL1Plugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code = FetchL1Plugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg = FetchL1Plugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid}}};
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2];
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[0] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 && (! 1'b0));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[1] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 && (! _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[2] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1})));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[3] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1}})));
  end

  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = (((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception}} : 39'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1}} : 39'h0)) | ((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2}} : 39'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3}} : 39'h0)));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[38 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = PrivilegedPlugin_logic_harts_0_m_status_mpp;
  assign TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b11;
  assign TrapPlugin_logic_harts_0_trap_exception_code = TrapPlugin_logic_harts_0_trap_pending_state_code;
  assign TrapPlugin_logic_harts_0_trap_exception_targetPrivilege = ((PrivilegedPlugin_logic_harts_0_privilege < TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped) ? TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_commitMask = {(((execute_ctrl5_down_LANE_SEL_lane1 && execute_ctrl5_down_isReady) && (! execute_lane1_ctrls_5_downIsCancel)) && execute_ctrl5_down_COMMIT_lane1),(((execute_ctrl5_down_LANE_SEL_lane0 && execute_ctrl5_down_isReady) && (! execute_lane0_ctrls_5_downIsCancel)) && execute_ctrl5_down_COMMIT_lane0)};
  assign TrapPlugin_logic_harts_0_trap_trigger_oh = {(((execute_ctrl4_down_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_downIsCancel)) && execute_ctrl4_down_TRAP_lane1),(((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_TRAP_lane0)};
  assign TrapPlugin_logic_harts_0_trap_trigger_valid = (|TrapPlugin_logic_harts_0_trap_trigger_oh);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_pc = TrapPlugin_logic_harts_0_trap_trigger_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 = TrapPlugin_logic_harts_0_trap_trigger_oh[1];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_interrupt = 1'bx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_interrupt = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_code = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_code = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_historyPort_payload_history = TrapPlugin_logic_harts_0_trap_pending_history;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_pcPort_payload_fault = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_pending_pc;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantExit = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
        TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantKill = 1'b0;
  assign TrapPlugin_logic_harts_0_trap_fsm_inflightTrap = (|{execute_lane1_logic_trapPending[0],{execute_lane0_logic_trapPending[0],{DispatchPlugin_logic_trapPendings[0],decode_logic_trapPending[0]}}});
  assign TrapPlugin_logic_harts_0_trap_fsm_holdPort = (TrapPlugin_logic_harts_0_trap_fsm_inflightTrap || (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING)));
  assign TrapPlugin_api_harts_0_fsmBusy = (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b1;
            end
            4'b0110 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt = ((TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0000) && TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege : TrapPlugin_logic_harts_0_trap_exception_targetPrivilege);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval = ((! TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt) ? TrapPlugin_logic_harts_0_trap_pending_state_tval : 32'h0);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code : TrapPlugin_logic_harts_0_trap_pending_state_code);
  assign TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0 = (! TrapPlugin_logic_initHold);
  assign TrapPlugin_logic_harts_0_trap_fsm_jumpOffset = ((|{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b1000),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0110),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0010),(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0101)}}}) ? TrapPlugin_logic_harts_0_trap_pending_slices : 2'b00);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak = 1'b0;
  assign when_TrapPlugin_l556 = (TrapPlugin_logic_harts_0_crsPorts_read_valid && TrapPlugin_logic_harts_0_crsPorts_read_ready);
  assign TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign PcPlugin_logic_forcedSpawn = (|{TrapPlugin_logic_harts_0_trap_pcPort_valid,{late1_BranchPlugin_logic_pcPort_valid,{early1_BranchPlugin_logic_pcPort_valid,{late0_BranchPlugin_logic_pcPort_valid,{early0_BranchPlugin_logic_pcPort_valid,BtbPlugin_logic_pcPort_valid}}}}});
  assign PcPlugin_logic_harts_0_self_pc = (PcPlugin_logic_harts_0_self_state + _zz_PcPlugin_logic_harts_0_self_pc);
  assign PcPlugin_logic_harts_0_self_flow_valid = 1'b1;
  assign PcPlugin_logic_harts_0_self_flow_payload_fault = PcPlugin_logic_harts_0_self_fault;
  assign PcPlugin_logic_harts_0_self_flow_payload_pc = PcPlugin_logic_harts_0_self_pc;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid = (&((! early1_BranchPlugin_logic_pcPort_valid) || (early0_BranchPlugin_logic_pcPort_payload_laneAge < early1_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid = (&((! late1_BranchPlugin_logic_pcPort_valid) || (late0_BranchPlugin_logic_pcPort_payload_laneAge < late1_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid = (&((! early0_BranchPlugin_logic_pcPort_valid) || (early1_BranchPlugin_logic_pcPort_payload_laneAge < early0_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid = (&((! late0_BranchPlugin_logic_pcPort_valid) || (late1_BranchPlugin_logic_pcPort_payload_laneAge < late0_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_valids_0 = ((TrapPlugin_logic_harts_0_trap_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_1 = ((late0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_2 = ((late1_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_3 = ((early0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_4 = ((early1_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_5 = ((BtbPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_6 = ((PcPlugin_logic_harts_0_self_flow_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid);
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh = {PcPlugin_logic_harts_0_aggregator_valids_6,{PcPlugin_logic_harts_0_aggregator_valids_5,{PcPlugin_logic_harts_0_aggregator_valids_4,{PcPlugin_logic_harts_0_aggregator_valids_3,{PcPlugin_logic_harts_0_aggregator_valids_2,{PcPlugin_logic_harts_0_aggregator_valids_1,PcPlugin_logic_harts_0_aggregator_valids_0}}}}}};
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_1 = _zz_PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_2 = _zz_PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_3 = _zz_PcPlugin_logic_harts_0_aggregator_oh[2];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_4 = _zz_PcPlugin_logic_harts_0_aggregator_oh[3];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_5 = _zz_PcPlugin_logic_harts_0_aggregator_oh[4];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_6 = _zz_PcPlugin_logic_harts_0_aggregator_oh[5];
  always @(*) begin
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[0] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[1] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_2 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_1));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[2] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_3 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[3] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_4 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[4] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_5 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_8));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[5] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_6 && (! (_zz_PcPlugin_logic_harts_0_aggregator_oh_5 || _zz_PcPlugin_logic_harts_0_aggregator_oh_8)));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[6] = (_zz_PcPlugin_logic_harts_0_aggregator_oh[6] && (! ((|{_zz_PcPlugin_logic_harts_0_aggregator_oh_6,_zz_PcPlugin_logic_harts_0_aggregator_oh_5}) || _zz_PcPlugin_logic_harts_0_aggregator_oh_8)));
  end

  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_8 = (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_4,{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}}});
  assign PcPlugin_logic_harts_0_aggregator_oh = _zz_PcPlugin_logic_harts_0_aggregator_oh_7;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target = PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_2 = PcPlugin_logic_harts_0_aggregator_oh[2];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_3 = PcPlugin_logic_harts_0_aggregator_oh[3];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_4 = PcPlugin_logic_harts_0_aggregator_oh[4];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_5 = PcPlugin_logic_harts_0_aggregator_oh[6];
  assign PcPlugin_logic_harts_0_aggregator_target = ((((_zz_PcPlugin_logic_harts_0_aggregator_target ? _zz_PcPlugin_logic_harts_0_aggregator_target_6 : _zz_PcPlugin_logic_harts_0_aggregator_target_7) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? _zz_PcPlugin_logic_harts_0_aggregator_target_8 : _zz_PcPlugin_logic_harts_0_aggregator_target_9)) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? _zz_PcPlugin_logic_harts_0_aggregator_target_10 : _zz_PcPlugin_logic_harts_0_aggregator_target_11) | (_zz_PcPlugin_logic_harts_0_aggregator_target_3 ? _zz_PcPlugin_logic_harts_0_aggregator_target_12 : _zz_PcPlugin_logic_harts_0_aggregator_target_13))) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_4 ? early1_BranchPlugin_logic_pcPort_payload_pc : 32'h0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_5 ? PcPlugin_logic_harts_0_self_flow_payload_pc : 32'h0)));
  assign PcPlugin_logic_harts_0_aggregator_fault = _zz_PcPlugin_logic_harts_0_aggregator_fault[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_oh[5];
  assign when_PcPlugin_l80 = (|_zz_PcPlugin_logic_harts_0_aggregator_fault_1);
  assign PcPlugin_logic_harts_0_holdComb = (|TrapPlugin_logic_harts_0_trap_fsm_holdPort);
  assign PcPlugin_logic_harts_0_output_valid = (! PcPlugin_logic_harts_0_holdReg);
  assign PcPlugin_logic_harts_0_output_payload_fault = PcPlugin_logic_harts_0_aggregator_fault_1;
  always @(*) begin
    PcPlugin_logic_harts_0_output_payload_pc = PcPlugin_logic_harts_0_aggregator_target_1;
    PcPlugin_logic_harts_0_output_payload_pc[0 : 0] = 1'b0;
  end

  assign PcPlugin_logic_harts_0_output_fire = (PcPlugin_logic_harts_0_output_valid && PcPlugin_logic_harts_0_output_ready);
  assign fetch_logic_ctrls_0_up_valid = PcPlugin_logic_harts_0_output_valid;
  assign PcPlugin_logic_harts_0_output_ready = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_0_up_Fetch_WORD_PC = PcPlugin_logic_harts_0_output_payload_pc;
  assign fetch_logic_ctrls_0_up_Fetch_PC_FAULT = PcPlugin_logic_harts_0_output_payload_fault;
  always @(*) begin
    fetch_logic_ctrls_0_up_Fetch_ID = 10'bxxxxxxxxxx;
    fetch_logic_ctrls_0_up_Fetch_ID = PcPlugin_logic_harts_0_self_id;
  end

  assign PcPlugin_logic_holdHalter_doIt = PcPlugin_logic_harts_0_holdComb;
  assign fetch_logic_ctrls_0_haltRequest_PcPlugin_l133 = PcPlugin_logic_holdHalter_doIt;
  assign CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_interface_fire = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_interface_fire = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_inject_csrAddress = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign CsrAccessPlugin_logic_fsm_inject_immZero = (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0);
  assign CsrAccessPlugin_logic_fsm_inject_srcZero = (execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 ? CsrAccessPlugin_logic_fsm_inject_immZero : (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0));
  assign CsrAccessPlugin_logic_fsm_inject_csrWrite = (! (execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 && CsrAccessPlugin_logic_fsm_inject_srcZero));
  assign CsrAccessPlugin_logic_fsm_inject_csrRead = (! ((! execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0) && (! execute_ctrl2_up_RD_ENABLE_lane0)));
  assign COMB_CSR_2047 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7ff);
  assign COMB_CSR_1952 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a0);
  assign COMB_CSR_1953 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a1);
  assign COMB_CSR_1954 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a2);
  assign COMB_CSR_3857 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf11);
  assign COMB_CSR_3858 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf12);
  assign COMB_CSR_3859 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf13);
  assign COMB_CSR_3860 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf14);
  assign COMB_CSR_769 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h301);
  assign COMB_CSR_768 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300);
  assign COMB_CSR_834 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h342);
  assign COMB_CSR_836 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h344);
  assign COMB_CSR_772 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h304);
  assign COMB_CSR_3 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h003);
  assign COMB_CSR_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h002);
  assign COMB_CSR_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h001);
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter = (|(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305));
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter = (|(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341));
  assign COMB_CSR_FpuCsrPlugin_logic_csrDirty = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h001),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h003),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h002)}});
  assign COMB_CSR_CsrRamPlugin_csrMapper_selFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h340),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h343),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)}}});
  assign COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h003),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h002),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300)}});
  assign CsrAccessPlugin_logic_fsm_inject_implemented = (|{COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter,{COMB_CSR_CsrRamPlugin_csrMapper_selFilter,{COMB_CSR_FpuCsrPlugin_logic_csrDirty,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter,{COMB_CSR_1,{COMB_CSR_2,{COMB_CSR_3,{COMB_CSR_772,{COMB_CSR_836,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_1}}}}}}}}}}});
  assign CsrAccessPlugin_logic_fsm_inject_onDecodeDo = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign when_CsrAccessPlugin_l155 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter);
  assign CsrAccessPlugin_logic_fsm_inject_trap = ((! CsrAccessPlugin_logic_fsm_inject_implemented) || CsrAccessPlugin_bus_decode_exception);
  assign CsrAccessPlugin_bus_decode_read = CsrAccessPlugin_logic_fsm_inject_csrRead;
  assign CsrAccessPlugin_bus_decode_write = CsrAccessPlugin_logic_fsm_inject_csrWrite;
  assign CsrAccessPlugin_bus_decode_address = CsrAccessPlugin_logic_fsm_inject_csrAddress;
  assign CsrAccessPlugin_logic_fsm_interface_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rs1 = execute_ctrl2_up_integer_RS1_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_uop = execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doImm = execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doMask = execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doClear = execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdEnable = execute_ctrl2_up_RD_ENABLE_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdPhys = execute_ctrl2_down_RD_PHYS_lane0;
  assign CsrAccessPlugin_logic_fsm_inject_freeze = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (! CsrAccessPlugin_logic_fsm_inject_unfreeze));
  always @(*) begin
    CsrAccessPlugin_logic_flushPort_valid = 1'b0;
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      CsrAccessPlugin_logic_flushPort_valid = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_flushPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_flushPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_trapPort_valid = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_trapPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_exception = 1'b1;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_exception = 1'b0;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_code = 4'b0010;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_code = CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_trapPort_payload_tval = execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_trapPort_payload_arg = 2'b00;
  assign CsrAccessPlugin_logic_trapPort_payload_laneAge = execute_ctrl2_down_LANE_AGE_lane0;
  assign when_CsrAccessPlugin_l197 = (! execute_freeze_valid);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = CsrAccessPlugin_logic_fsm_interface_read;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l296) begin
          CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = CsrAccessPlugin_logic_fsm_interface_read;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_read_valid = CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  assign CsrAccessPlugin_bus_read_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  assign CsrAccessPlugin_bus_read_moving = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l252 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30)))) | ((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46))) | (CsrRamPlugin_csrMapper_withRead ? CsrRamPlugin_csrMapper_read_data : 32'h0)));
  assign CsrAccessPlugin_bus_read_data = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  assign CsrAccessPlugin_bus_read_toWriteBits = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = REG_CSR_3;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue = 1'b1;
  assign CsrAccessPlugin_bus_write_moving = (! CsrAccessPlugin_bus_write_halt);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (CsrAccessPlugin_logic_fsm_interface_doImm ? _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : CsrAccessPlugin_logic_fsm_interface_rs1);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (CsrAccessPlugin_logic_fsm_interface_doClear ? (CsrAccessPlugin_logic_fsm_interface_aluInput & (~ CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (CsrAccessPlugin_logic_fsm_interface_aluInput | CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (CsrAccessPlugin_logic_fsm_interface_doMask ? CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  always @(*) begin
    CsrAccessPlugin_bus_write_bits = CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l343) begin
      CsrAccessPlugin_bus_write_bits[1 : 0] = 2'b00;
    end
    if(when_CsrAccessPlugin_l343_1) begin
      CsrAccessPlugin_bus_write_bits[0 : 0] = 1'b0;
    end
  end

  assign CsrAccessPlugin_bus_write_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = CsrAccessPlugin_logic_fsm_interface_write;
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l325) begin
          CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = CsrAccessPlugin_logic_fsm_interface_write;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_write_valid = CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  assign when_CsrAccessPlugin_l346 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_2047);
  assign when_CsrAccessPlugin_l346_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign when_CsrAccessPlugin_l346_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l346_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l346_4 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_3);
  assign _zz_FpuCsrPlugin_api_flags_NX = CsrAccessPlugin_bus_write_bits[4 : 0];
  assign when_CsrAccessPlugin_l346_5 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_2);
  assign when_CsrAccessPlugin_l346_6 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_1);
  assign _zz_FpuCsrPlugin_api_flags_NX_1 = CsrAccessPlugin_bus_write_bits[4 : 0];
  assign when_CsrAccessPlugin_l343 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter);
  assign when_CsrAccessPlugin_l343_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter);
  assign when_CsrAccessPlugin_l346_7 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_FpuCsrPlugin_logic_csrDirty);
  assign when_CsrAccessPlugin_l343_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign CsrAccessPlugin_logic_wbWi_valid = execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  assign CsrAccessPlugin_logic_wbWi_payload = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign fetch_logic_ctrls_1_down_MMU_REFILL = 1'b0;
  assign fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
  assign fetch_logic_ctrls_1_down_MMU_TRANSLATED = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  assign fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = 1'b1;
  assign fetch_logic_ctrls_1_down_MMU_ALLOW_READ = 1'b1;
  assign fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = 1'b1;
  assign fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = 1'b0;
  assign fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
  assign fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION = 1'b1;
  assign execute_ctrl3_down_MMU_REFILL_lane0 = 1'b0;
  assign execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
  assign execute_ctrl3_down_MMU_TRANSLATED_lane0 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = 1'b1;
  assign execute_ctrl3_down_MMU_ALLOW_READ_lane0 = 1'b1;
  assign execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = 1'b1;
  assign execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = 1'b0;
  assign execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
  assign execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0 = 1'b1;
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(HistoryPlugin_logic_onFetch_ports_0_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_0_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_1_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_1_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_2_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_2_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_3_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_3_payload_history;
    end
  end

  assign HistoryPlugin_logic_onFetch_ports_0_valid = (|BtbPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_0_payload_history = BtbPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_1_valid = (|{early1_BranchPlugin_logic_historyPort_valid,early0_BranchPlugin_logic_historyPort_valid});
  assign _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history = (((early0_BranchPlugin_logic_historyPort_valid && (&(! (early1_BranchPlugin_logic_historyPort_valid && (early1_BranchPlugin_logic_historyPort_payload_age < early0_BranchPlugin_logic_historyPort_payload_age))))) ? {early0_BranchPlugin_logic_historyPort_payload_age,early0_BranchPlugin_logic_historyPort_payload_history} : 13'h0) | ((early1_BranchPlugin_logic_historyPort_valid && (&(! (early0_BranchPlugin_logic_historyPort_valid && (early0_BranchPlugin_logic_historyPort_payload_age < early1_BranchPlugin_logic_historyPort_payload_age))))) ? {early1_BranchPlugin_logic_historyPort_payload_age,early1_BranchPlugin_logic_historyPort_payload_history} : 13'h0));
  assign HistoryPlugin_logic_onFetch_ports_1_payload_history = _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history[11 : 0];
  assign HistoryPlugin_logic_onFetch_ports_1_payload_age = _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history[12 : 12];
  assign HistoryPlugin_logic_onFetch_ports_2_valid = (|{late1_BranchPlugin_logic_historyPort_valid,late0_BranchPlugin_logic_historyPort_valid});
  assign _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history = (((late0_BranchPlugin_logic_historyPort_valid && (&(! (late1_BranchPlugin_logic_historyPort_valid && (late1_BranchPlugin_logic_historyPort_payload_age < late0_BranchPlugin_logic_historyPort_payload_age))))) ? {late0_BranchPlugin_logic_historyPort_payload_age,late0_BranchPlugin_logic_historyPort_payload_history} : 13'h0) | ((late1_BranchPlugin_logic_historyPort_valid && (&(! (late0_BranchPlugin_logic_historyPort_valid && (late0_BranchPlugin_logic_historyPort_payload_age < late1_BranchPlugin_logic_historyPort_payload_age))))) ? {late1_BranchPlugin_logic_historyPort_payload_age,late1_BranchPlugin_logic_historyPort_payload_history} : 13'h0));
  assign HistoryPlugin_logic_onFetch_ports_2_payload_history = _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history[11 : 0];
  assign HistoryPlugin_logic_onFetch_ports_2_payload_age = _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history[12 : 12];
  assign HistoryPlugin_logic_onFetch_ports_3_valid = (|TrapPlugin_logic_harts_0_trap_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_3_payload_history = TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  assign fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{CsrRamPlugin_csrMapper_write_valid,TrapPlugin_logic_harts_0_crsPorts_write_valid}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign _zz_CsrRamPlugin_csrMapper_write_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = (((_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_address : 2'b00) | (_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_address : 2'b00)) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_address : 2'b00));
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = (((_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_data : 32'h0) | (_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_data : 32'h0)) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_data : 32'h0));
  assign TrapPlugin_logic_harts_0_crsPorts_write_ready = _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  assign CsrRamPlugin_csrMapper_write_ready = _zz_CsrRamPlugin_csrMapper_write_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {CsrRamPlugin_csrMapper_read_valid,TrapPlugin_logic_harts_0_crsPorts_read_valid};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_CsrRamPlugin_logic_readLogic_sel = CsrRamPlugin_logic_readLogic_oh[1];
  assign CsrRamPlugin_logic_readLogic_sel = _zz_CsrRamPlugin_logic_readLogic_sel;
  assign CsrRamPlugin_logic_readLogic_port_rsp = CsrRamPlugin_logic_mem_spinal_port1;
  assign CsrRamPlugin_logic_readLogic_port_cmd_valid = (((|CsrRamPlugin_logic_readLogic_oh) && (! CsrRamPlugin_logic_writeLogic_port_valid)) && (! CsrRamPlugin_logic_readLogic_busy));
  assign CsrRamPlugin_logic_readLogic_port_cmd_payload = _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  assign TrapPlugin_logic_harts_0_crsPorts_read_ready = CsrRamPlugin_logic_readLogic_ohReg[0];
  assign CsrRamPlugin_csrMapper_read_ready = CsrRamPlugin_logic_readLogic_ohReg[1];
  assign TrapPlugin_logic_harts_0_crsPorts_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_csrMapper_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[2];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[1:0];
  assign CsrRamPlugin_setup_initPort_data = 32'h0;
  assign execute_lane0_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS1_port_address = execute_ctrl0_down_RS1_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_integer_RS1_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl2_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[1] = (((execute_ctrl2_up_LANE_SEL_lane1 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl2_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[2] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[3] = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[4] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[5] = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[6] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[7] = (((execute_ctrl5_up_LANE_SEL_lane1 && execute_ctrl5_up_RD_ENABLE_lane1) && (execute_ctrl5_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_integer_RS1_bypassEnables[8] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS1_bypassEnables;
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[4];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[5];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[6];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[7];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS1_sel[0] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[1] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[2] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS1_sel[3] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS1_sel[4] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3));
    _zz_execute_lane0_bypasser_integer_RS1_sel[5] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5 && (! (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 || execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS1_sel[6] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6 && (! (execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5 || execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS1_sel[7] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7 && (! (execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6 || execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS1_sel[8] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8 && (! (execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7 || execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
  end

  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4}});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4}}});
  assign execute_lane0_bypasser_integer_RS1_sel = _zz_execute_lane0_bypasser_integer_RS1_sel;
  assign _zz_execute_ctrl1_down_integer_RS1_lane0 = execute_lane0_bypasser_integer_RS1_sel[8 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS1_lane0_1 = ((((_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1 ? execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_1) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_2 ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_3)) | ((_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_4 ? execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_5) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_6 ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_7))) | (((_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_8 ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_9) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_10 ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_11)) | ((_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_12 ? execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_13) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_14 ? execute_lane0_bypasser_integer_RS1_port_data : _zz__zz_execute_ctrl1_down_integer_RS1_lane0_1_15))));
    if(when_ExecuteLanePlugin_l196) begin
      _zz_execute_ctrl1_down_integer_RS1_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS1_lane0 = _zz_execute_ctrl1_down_integer_RS1_lane0_1;
  assign when_ExecuteLanePlugin_l196 = execute_lane0_bypasser_integer_RS1_sel[0];
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit = (execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit && (! (|{execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1,execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0})));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit = (execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit = (execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit && (! (|{execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1,execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0})));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits = {execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit,{execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit,execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit}};
  assign _zz_execute_ctrl2_integer_RS1_lane0_bypass = {execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits,(! (|execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits))};
  assign execute_ctrl2_integer_RS1_lane0_bypass = (((_zz_execute_ctrl2_integer_RS1_lane0_bypass[0] ? execute_ctrl2_up_integer_RS1_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS1_lane0_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl2_integer_RS1_lane0_bypass[2] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS1_lane0_bypass[3] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0)));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl3_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl3_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit = (execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl3_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl3_down_RS1_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit = (execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits = {execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit,execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit};
  assign _zz_execute_ctrl3_integer_RS1_lane0_bypass = {execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits,(! (|execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits))};
  assign execute_ctrl3_integer_RS1_lane0_bypass = (((_zz_execute_ctrl3_integer_RS1_lane0_bypass[0] ? execute_ctrl3_up_integer_RS1_lane0 : 32'h0) | (_zz_execute_ctrl3_integer_RS1_lane0_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_execute_ctrl3_integer_RS1_lane0_bypass[2] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane0_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS2_port_address = execute_ctrl0_down_RS2_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_integer_RS2_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl2_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[1] = (((execute_ctrl2_up_LANE_SEL_lane1 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl2_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[2] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[3] = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[4] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[5] = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[6] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[7] = (((execute_ctrl5_up_LANE_SEL_lane1 && execute_ctrl5_up_RD_ENABLE_lane1) && (execute_ctrl5_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_integer_RS2_bypassEnables[8] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS2_bypassEnables;
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[4];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[5];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[6];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[7];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS2_sel[0] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[1] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[2] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS2_sel[3] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS2_sel[4] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3));
    _zz_execute_lane0_bypasser_integer_RS2_sel[5] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5 && (! (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 || execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS2_sel[6] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6 && (! (execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5 || execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS2_sel[7] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7 && (! (execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6 || execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_integer_RS2_sel[8] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8 && (! (execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7 || execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
  end

  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4}});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4}}});
  assign execute_lane0_bypasser_integer_RS2_sel = _zz_execute_lane0_bypasser_integer_RS2_sel;
  assign _zz_execute_ctrl1_down_integer_RS2_lane0 = execute_lane0_bypasser_integer_RS2_sel[8 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS2_lane0_1 = ((((_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1 ? execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_1) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_2 ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_3)) | ((_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_4 ? execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_5) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_6 ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_7))) | (((_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_8 ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_9) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_10 ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_11)) | ((_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_12 ? execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_13) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_14 ? execute_lane0_bypasser_integer_RS2_port_data : _zz__zz_execute_ctrl1_down_integer_RS2_lane0_1_15))));
    if(when_ExecuteLanePlugin_l196_1) begin
      _zz_execute_ctrl1_down_integer_RS2_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS2_lane0 = _zz_execute_ctrl1_down_integer_RS2_lane0_1;
  assign when_ExecuteLanePlugin_l196_1 = execute_lane0_bypasser_integer_RS2_sel[0];
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit = (execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit && (! (|{execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1,execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0})));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit = (execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane0)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit = (execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit && (! (|{execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1,execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0})));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits = {execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit,{execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit,execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit}};
  assign _zz_execute_ctrl2_integer_RS2_lane0_bypass = {execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits,(! (|execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits))};
  assign execute_ctrl2_integer_RS2_lane0_bypass = (((_zz_execute_ctrl2_integer_RS2_lane0_bypass[0] ? execute_ctrl2_up_integer_RS2_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS2_lane0_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl2_integer_RS2_lane0_bypass[2] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS2_lane0_bypass[3] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0)));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl3_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl3_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit = (execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl3_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl3_down_RS2_RFID_lane0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit = (execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits = {execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit,execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit};
  assign _zz_execute_ctrl3_integer_RS2_lane0_bypass = {execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits,(! (|execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits))};
  assign execute_ctrl3_integer_RS2_lane0_bypass = (((_zz_execute_ctrl3_integer_RS2_lane0_bypass[0] ? execute_ctrl3_up_integer_RS2_lane0 : 32'h0) | (_zz_execute_ctrl3_integer_RS2_lane0_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_execute_ctrl3_integer_RS2_lane0_bypass[2] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane0_bypasser_float_RS1_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_float_RS1_port_address = execute_ctrl0_down_RS1_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_float_RS1_bypassEnables[0] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[1] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[2] = (((execute_ctrl6_up_LANE_SEL_lane0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl6_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[3] = (((execute_ctrl7_up_LANE_SEL_lane0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl7_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[4] = (((execute_ctrl8_up_LANE_SEL_lane0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl8_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[5] = (((execute_ctrl9_up_LANE_SEL_lane0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl9_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[6] = (((execute_ctrl10_up_LANE_SEL_lane0 && execute_ctrl10_up_RD_ENABLE_lane0) && (execute_ctrl10_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl10_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[7] = (((execute_ctrl11_up_LANE_SEL_lane0 && execute_ctrl11_up_RD_ENABLE_lane0) && (execute_ctrl11_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl11_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[8] = (((execute_ctrl12_up_LANE_SEL_lane0 && execute_ctrl12_up_RD_ENABLE_lane0) && (execute_ctrl12_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && (execute_ctrl12_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane0));
    execute_lane0_bypasser_float_RS1_bypassEnables[9] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0 = execute_lane0_bypasser_float_RS1_bypassEnables;
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[4];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_5 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[5];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_6 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[6];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_7 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[7];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_8 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[8];
  assign execute_lane0_bypasser_float_RS1_bypassEnables_bools_9 = _zz_execute_lane0_bypasser_float_RS1_bypassEnables_bools_0[9];
  always @(*) begin
    _zz_execute_lane0_bypasser_float_RS1_sel[0] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_float_RS1_sel[1] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_1 && (! execute_lane0_bypasser_float_RS1_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_float_RS1_sel[2] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_2 && (! execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_float_RS1_sel[3] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_3 && (! execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_float_RS1_sel[4] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_4 && (! execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3));
    _zz_execute_lane0_bypasser_float_RS1_sel[5] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_5 && (! (execute_lane0_bypasser_float_RS1_bypassEnables_bools_4 || execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS1_sel[6] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_6 && (! (execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_5 || execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS1_sel[7] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_7 && (! (execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_6 || execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS1_sel[8] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_8 && (! (execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_7 || execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS1_sel[9] = (execute_lane0_bypasser_float_RS1_bypassEnables_bools_9 && (! (execute_lane0_bypasser_float_RS1_bypassEnables_bools_8 || execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_7)));
  end

  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_1,execute_lane0_bypasser_float_RS1_bypassEnables_bools_0});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_1,execute_lane0_bypasser_float_RS1_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_3,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_1,execute_lane0_bypasser_float_RS1_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_5 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_5,execute_lane0_bypasser_float_RS1_bypassEnables_bools_4});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_6 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_5,execute_lane0_bypasser_float_RS1_bypassEnables_bools_4}});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_7 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_bools_7,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS1_bypassEnables_bools_5,execute_lane0_bypasser_float_RS1_bypassEnables_bools_4}}});
  assign execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_7 = (|{execute_lane0_bypasser_float_RS1_bypassEnables_range_4_to_7,execute_lane0_bypasser_float_RS1_bypassEnables_range_0_to_3});
  assign execute_lane0_bypasser_float_RS1_sel = _zz_execute_lane0_bypasser_float_RS1_sel;
  assign execute_ctrl1_down_float_RS1_lane0 = (((((_zz_execute_ctrl1_down_float_RS1_lane0 ? execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_1) | (_zz_execute_ctrl1_down_float_RS1_lane0_2 ? execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_3)) | ((_zz_execute_ctrl1_down_float_RS1_lane0_4 ? execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_5) | (_zz_execute_ctrl1_down_float_RS1_lane0_6 ? execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_7))) | (((_zz_execute_ctrl1_down_float_RS1_lane0_8 ? execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_9) | (_zz_execute_ctrl1_down_float_RS1_lane0_10 ? execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_11)) | ((_zz_execute_ctrl1_down_float_RS1_lane0_12 ? execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_13) | (_zz_execute_ctrl1_down_float_RS1_lane0_14 ? execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS1_lane0_15)))) | ((execute_lane0_bypasser_float_RS1_sel[8] ? execute_ctrl12_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (execute_lane0_bypasser_float_RS1_sel[9] ? execute_lane0_bypasser_float_RS1_port_data : 64'h0)));
  assign execute_lane0_bypasser_float_RS2_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_float_RS2_port_address = execute_ctrl0_down_RS2_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_float_RS2_bypassEnables[0] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[1] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[2] = (((execute_ctrl6_up_LANE_SEL_lane0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl6_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[3] = (((execute_ctrl7_up_LANE_SEL_lane0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl7_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[4] = (((execute_ctrl8_up_LANE_SEL_lane0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl8_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[5] = (((execute_ctrl9_up_LANE_SEL_lane0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl9_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[6] = (((execute_ctrl10_up_LANE_SEL_lane0 && execute_ctrl10_up_RD_ENABLE_lane0) && (execute_ctrl10_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl10_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[7] = (((execute_ctrl11_up_LANE_SEL_lane0 && execute_ctrl11_up_RD_ENABLE_lane0) && (execute_ctrl11_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl11_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[8] = (((execute_ctrl12_up_LANE_SEL_lane0 && execute_ctrl12_up_RD_ENABLE_lane0) && (execute_ctrl12_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && (execute_ctrl12_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane0));
    execute_lane0_bypasser_float_RS2_bypassEnables[9] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0 = execute_lane0_bypasser_float_RS2_bypassEnables;
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[4];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_5 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[5];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_6 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[6];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_7 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[7];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_8 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[8];
  assign execute_lane0_bypasser_float_RS2_bypassEnables_bools_9 = _zz_execute_lane0_bypasser_float_RS2_bypassEnables_bools_0[9];
  always @(*) begin
    _zz_execute_lane0_bypasser_float_RS2_sel[0] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_float_RS2_sel[1] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_1 && (! execute_lane0_bypasser_float_RS2_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_float_RS2_sel[2] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_2 && (! execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_float_RS2_sel[3] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_3 && (! execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_float_RS2_sel[4] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_4 && (! execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3));
    _zz_execute_lane0_bypasser_float_RS2_sel[5] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_5 && (! (execute_lane0_bypasser_float_RS2_bypassEnables_bools_4 || execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS2_sel[6] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_6 && (! (execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_5 || execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS2_sel[7] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_7 && (! (execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_6 || execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS2_sel[8] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_8 && (! (execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_7 || execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS2_sel[9] = (execute_lane0_bypasser_float_RS2_bypassEnables_bools_9 && (! (execute_lane0_bypasser_float_RS2_bypassEnables_bools_8 || execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_7)));
  end

  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_1,execute_lane0_bypasser_float_RS2_bypassEnables_bools_0});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_1,execute_lane0_bypasser_float_RS2_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_3,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_1,execute_lane0_bypasser_float_RS2_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_5 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_5,execute_lane0_bypasser_float_RS2_bypassEnables_bools_4});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_6 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_5,execute_lane0_bypasser_float_RS2_bypassEnables_bools_4}});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_7 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_bools_7,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS2_bypassEnables_bools_5,execute_lane0_bypasser_float_RS2_bypassEnables_bools_4}}});
  assign execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_7 = (|{execute_lane0_bypasser_float_RS2_bypassEnables_range_4_to_7,execute_lane0_bypasser_float_RS2_bypassEnables_range_0_to_3});
  assign execute_lane0_bypasser_float_RS2_sel = _zz_execute_lane0_bypasser_float_RS2_sel;
  assign execute_ctrl1_down_float_RS2_lane0 = (((((_zz_execute_ctrl1_down_float_RS2_lane0 ? execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_1) | (_zz_execute_ctrl1_down_float_RS2_lane0_2 ? execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_3)) | ((_zz_execute_ctrl1_down_float_RS2_lane0_4 ? execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_5) | (_zz_execute_ctrl1_down_float_RS2_lane0_6 ? execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_7))) | (((_zz_execute_ctrl1_down_float_RS2_lane0_8 ? execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_9) | (_zz_execute_ctrl1_down_float_RS2_lane0_10 ? execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_11)) | ((_zz_execute_ctrl1_down_float_RS2_lane0_12 ? execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_13) | (_zz_execute_ctrl1_down_float_RS2_lane0_14 ? execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS2_lane0_15)))) | ((execute_lane0_bypasser_float_RS2_sel[8] ? execute_ctrl12_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (execute_lane0_bypasser_float_RS2_sel[9] ? execute_lane0_bypasser_float_RS2_port_data : 64'h0)));
  assign execute_lane0_bypasser_float_RS3_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_float_RS3_port_address = execute_ctrl0_down_RS3_PHYS_lane0[4 : 0];
  always @(*) begin
    execute_lane0_bypasser_float_RS3_bypassEnables[0] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[1] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[2] = (((execute_ctrl6_up_LANE_SEL_lane0 && execute_ctrl6_up_RD_ENABLE_lane0) && (execute_ctrl6_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl6_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[3] = (((execute_ctrl7_up_LANE_SEL_lane0 && execute_ctrl7_up_RD_ENABLE_lane0) && (execute_ctrl7_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl7_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[4] = (((execute_ctrl8_up_LANE_SEL_lane0 && execute_ctrl8_up_RD_ENABLE_lane0) && (execute_ctrl8_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl8_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[5] = (((execute_ctrl9_up_LANE_SEL_lane0 && execute_ctrl9_up_RD_ENABLE_lane0) && (execute_ctrl9_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl9_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[6] = (((execute_ctrl10_up_LANE_SEL_lane0 && execute_ctrl10_up_RD_ENABLE_lane0) && (execute_ctrl10_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl10_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[7] = (((execute_ctrl11_up_LANE_SEL_lane0 && execute_ctrl11_up_RD_ENABLE_lane0) && (execute_ctrl11_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl11_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[8] = (((execute_ctrl12_up_LANE_SEL_lane0 && execute_ctrl12_up_RD_ENABLE_lane0) && (execute_ctrl12_down_RD_PHYS_lane0 == execute_ctrl1_down_RS3_PHYS_lane0)) && (execute_ctrl12_down_RD_RFID_lane0 == execute_ctrl1_down_RS3_RFID_lane0));
    execute_lane0_bypasser_float_RS3_bypassEnables[9] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0 = execute_lane0_bypasser_float_RS3_bypassEnables;
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[4];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_5 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[5];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_6 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[6];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_7 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[7];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_8 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[8];
  assign execute_lane0_bypasser_float_RS3_bypassEnables_bools_9 = _zz_execute_lane0_bypasser_float_RS3_bypassEnables_bools_0[9];
  always @(*) begin
    _zz_execute_lane0_bypasser_float_RS3_sel[0] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_float_RS3_sel[1] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_1 && (! execute_lane0_bypasser_float_RS3_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_float_RS3_sel[2] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_2 && (! execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_float_RS3_sel[3] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_3 && (! execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_float_RS3_sel[4] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_4 && (! execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3));
    _zz_execute_lane0_bypasser_float_RS3_sel[5] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_5 && (! (execute_lane0_bypasser_float_RS3_bypassEnables_bools_4 || execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS3_sel[6] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_6 && (! (execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_5 || execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS3_sel[7] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_7 && (! (execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_6 || execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS3_sel[8] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_8 && (! (execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_7 || execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3)));
    _zz_execute_lane0_bypasser_float_RS3_sel[9] = (execute_lane0_bypasser_float_RS3_bypassEnables_bools_9 && (! (execute_lane0_bypasser_float_RS3_bypassEnables_bools_8 || execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_7)));
  end

  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_1,execute_lane0_bypasser_float_RS3_bypassEnables_bools_0});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_1,execute_lane0_bypasser_float_RS3_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_3,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_2,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_1,execute_lane0_bypasser_float_RS3_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_5 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_5,execute_lane0_bypasser_float_RS3_bypassEnables_bools_4});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_6 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_5,execute_lane0_bypasser_float_RS3_bypassEnables_bools_4}});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_7 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_bools_7,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_6,{execute_lane0_bypasser_float_RS3_bypassEnables_bools_5,execute_lane0_bypasser_float_RS3_bypassEnables_bools_4}}});
  assign execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_7 = (|{execute_lane0_bypasser_float_RS3_bypassEnables_range_4_to_7,execute_lane0_bypasser_float_RS3_bypassEnables_range_0_to_3});
  assign execute_lane0_bypasser_float_RS3_sel = _zz_execute_lane0_bypasser_float_RS3_sel;
  assign execute_ctrl1_down_float_RS3_lane0 = (((((_zz_execute_ctrl1_down_float_RS3_lane0 ? execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_1) | (_zz_execute_ctrl1_down_float_RS3_lane0_2 ? execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_3)) | ((_zz_execute_ctrl1_down_float_RS3_lane0_4 ? execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_5) | (_zz_execute_ctrl1_down_float_RS3_lane0_6 ? execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_7))) | (((_zz_execute_ctrl1_down_float_RS3_lane0_8 ? execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_9) | (_zz_execute_ctrl1_down_float_RS3_lane0_10 ? execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_11)) | ((_zz_execute_ctrl1_down_float_RS3_lane0_12 ? execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_13) | (_zz_execute_ctrl1_down_float_RS3_lane0_14 ? execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : _zz_execute_ctrl1_down_float_RS3_lane0_15)))) | ((execute_lane0_bypasser_float_RS3_sel[8] ? execute_ctrl12_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 : 64'h0) | (execute_lane0_bypasser_float_RS3_sel[9] ? execute_lane0_bypasser_float_RS3_port_data : 64'h0)));
  assign execute_lane0_logic_completions_onCtrl_0_port_valid = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_trap = execute_ctrl4_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_commit = execute_ctrl4_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_valid = (((execute_ctrl7_down_LANE_SEL_lane0 && execute_ctrl7_down_isReady) && (! execute_lane0_ctrls_7_downIsCancel)) && execute_ctrl7_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_uopId = execute_ctrl7_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_trap = execute_ctrl7_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_commit = execute_ctrl7_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_valid = (((execute_ctrl11_down_LANE_SEL_lane0 && execute_ctrl11_down_isReady) && (! execute_lane0_ctrls_11_downIsCancel)) && execute_ctrl11_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_uopId = execute_ctrl11_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_trap = execute_ctrl11_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_commit = execute_ctrl11_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_3_port_valid = (((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && execute_ctrl3_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_3_port_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_3_port_payload_trap = execute_ctrl3_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_3_port_payload_commit = execute_ctrl3_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_4_port_valid = (((execute_ctrl5_down_LANE_SEL_lane0 && execute_ctrl5_down_isReady) && (! execute_lane0_ctrls_5_downIsCancel)) && execute_ctrl5_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_4_port_payload_uopId = execute_ctrl5_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_4_port_payload_trap = execute_ctrl5_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_4_port_payload_commit = execute_ctrl5_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_5_port_valid = (((execute_ctrl8_down_LANE_SEL_lane0 && execute_ctrl8_down_isReady) && (! execute_lane0_ctrls_8_downIsCancel)) && execute_ctrl8_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_5_port_payload_uopId = execute_ctrl8_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_5_port_payload_trap = execute_ctrl8_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_5_port_payload_commit = execute_ctrl8_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_6_port_valid = (((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && execute_ctrl2_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_6_port_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_6_port_payload_trap = execute_ctrl2_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_6_port_payload_commit = execute_ctrl2_down_COMMIT_lane0;
  assign execute_lane0_logic_decoding_decodingBits = {execute_ctrl1_down_lane0_LAYER_SEL_lane0,execute_ctrl1_down_Decode_UOP_lane0};
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h100106060) == 33'h100006000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h100003064) == 33'h100003000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h100806060) == 33'h100806000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h101006060) == 33'h101006000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_4 = ((execute_lane0_logic_decoding_decodingBits & 33'h1000060e0) == 33'h100006080);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_5 = ((execute_lane0_logic_decoding_decodingBits & 33'h100006860) == 33'h100006800);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_6 = ((execute_lane0_logic_decoding_decodingBits & 33'h100406060) == 33'h100406000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_7 = ((execute_lane0_logic_decoding_decodingBits & 33'h100006260) == 33'h100006200);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_8 = ((execute_lane0_logic_decoding_decodingBits & 33'h100006460) == 33'h100006400);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_9 = ((execute_lane0_logic_decoding_decodingBits & 33'h100006160) == 33'h100006100);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000014) == 33'h100000014);
  always @(*) begin
    execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_10 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000070) == 33'h100000060);
  always @(*) begin
    execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h002004064) == 33'h002004020);
  always @(*) begin
    execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_11 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001048) == 33'h000001008);
  always @(*) begin
    execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000010) == 33'h0);
  always @(*) begin
    execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002070) == 33'h000002070);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001070) == 33'h000001070);
  always @(*) begin
    execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h00000003c) == 33'h000000004);
  assign _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h080000060) == 33'h000000040);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000070) == 33'h000000040);
  assign _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h010000060) == 33'h010000040);
  always @(*) begin
    execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0 = _zz_execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuClassPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuClassPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuClassPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuF2iPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuF2iPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuF2iPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0 = _zz_execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0 = _zz_execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h001d07fe4) == 33'h000106000);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000058) == 33'h0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001050) == 33'h0);
  always @(*) begin
    execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_AguPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h070000070) == 33'h000000050);
  always @(*) begin
    execute_ctrl1_down_FpuAddPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuAddPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuAddPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuMulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuMulPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h0d0000070) == 33'h040000050);
  always @(*) begin
    execute_ctrl1_down_FpuXxPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuXxPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuXxPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuDivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_FpuDivPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuDivPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0 = _zz_execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000014) == 33'h000000014);
  always @(*) begin
    execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h098000070) == 33'h010000050);
  always @(*) begin
    execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_5_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_3_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_6_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0 = _zz_execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_FpuFlagsWritebackPlugin_SEL_9_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0 = _zz_execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0_3[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h002004064) == 33'h002000020);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4 = ((execute_lane0_logic_decoding_decodingBits & 33'h0a0000070) == 33'h080000050);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5 = ((execute_lane0_logic_decoding_decodingBits & 33'h018000070) == 33'h018000050);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6 = ((execute_lane0_logic_decoding_decodingBits & 33'h050000070) == 33'h050000050);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000000) == 33'h0);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_4_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_7_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_7_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_7_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_11_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_11_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_11_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h030000050) == 33'h020000050);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_3_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_5_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_5_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_5_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_8_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_8_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_8_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_12 = ((execute_lane0_logic_decoding_decodingBits & 33'h100002070) == 33'h100000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_13 = ((execute_lane0_logic_decoding_decodingBits & 33'h100004070) == 33'h100000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_14 = ((execute_lane0_logic_decoding_decodingBits & 33'h102000070) == 33'h100000030);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_15 = ((execute_lane0_logic_decoding_decodingBits & 33'h100003060) == 33'h100000060);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_2_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0_4[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0_16[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000006000) == 33'h0);
  assign _zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000004) == 33'h000000004);
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000006004) == 33'h000002000);
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000003000) == 33'h000002000);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000004000) == 33'h0);
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001000) == 33'h000001000);
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = {(|{_zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0,{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0}})};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0[0];
  assign _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000008) == 33'h000000008);
  assign execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0[0];
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0);
  assign _zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000024) == 33'h0);
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000000070) == 33'h000000020),((execute_lane0_logic_decoding_decodingBits & 33'h001d07fa0) == 33'h000106000)}}),(|{((execute_lane0_logic_decoding_decodingBits & 33'h000000050) == 33'h0),_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1})};
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h010000020) == 33'h000000020);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000010) == 33'h000000010);
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = {(|{_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000002020) == 33'h000002000),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h008002000) == 33'h000002000)}}}),(|((execute_lane0_logic_decoding_decodingBits & 33'h000001010) == 33'h000001000))};
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000070) == 33'h100000010);
  assign execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_3_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h018000010) == 33'h018000010);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h020000010) == 33'h020000010);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000040) == 33'h0);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000020) == 33'h000000020);
  assign execute_ctrl1_down_BYPASSED_AT_4_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_4_lane0[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h040000010) == 33'h040000010);
  assign execute_ctrl1_down_BYPASSED_AT_5_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_5_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_6_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_6_lane0_1[0];
  assign execute_ctrl1_down_BYPASSED_AT_7_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_7_lane0_2[0];
  assign execute_ctrl1_down_BYPASSED_AT_8_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_8_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_9_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_9_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_10_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_3[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002050) == 33'h000002000);
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1[0];
  assign execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0[0];
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h00000000c) == 33'h000000004);
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1 = {(|_zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0),(|_zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0)};
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002000) == 33'h000002000);
  assign execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0[0];
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h080001000) == 33'h0);
  assign execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0[0];
  assign execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0[0];
  assign _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h012000000) == 33'h012000000),{((execute_lane0_logic_decoding_decodingBits & 33'h082000000) == 33'h082000000),{((execute_lane0_logic_decoding_decodingBits & 33'h002000010) == 33'h002000000),{((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1) == 33'h002000000),((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1_1) == 33'h040000010)}}}});
  assign _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0 = _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_1;
  assign _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2 = _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0;
  assign execute_ctrl1_down_FpuUtils_FORMAT_lane0 = _zz_execute_ctrl1_down_FpuUtils_FORMAT_lane0_2;
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h008000000) == 33'h0));
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_1;
  assign _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2 = _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0;
  assign execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0_2;
  assign execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0_1[0];
  assign execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0_1[0];
  assign execute_ctrl1_down_FpuCmpPlugin_LESS_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_LESS_lane0_1[0];
  assign execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0 = _zz_execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0[0];
  assign execute_ctrl1_down_AguPlugin_LOAD_lane0 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0[0];
  assign execute_ctrl1_down_AguPlugin_STORE_lane0 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0[0];
  assign execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0[0];
  assign execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0[0];
  assign execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1 = {(|((execute_lane0_logic_decoding_decodingBits & 33'h030001000) == 33'h010000000)),{(|{((execute_lane0_logic_decoding_decodingBits & 33'h020000000) == 33'h020000000),_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1}),(|{((execute_lane0_logic_decoding_decodingBits & 33'h000100000) == 33'h000100000),_zz_execute_ctrl1_down_BYPASSED_AT_10_lane0_1})}};
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  assign execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  assign execute_ctrl1_down_FpuAddPlugin_SUB_lane0 = _zz_execute_ctrl1_down_FpuAddPlugin_SUB_lane0[0];
  assign execute_ctrl1_down_FpuMulPlugin_FMA_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_FMA_lane0[0];
  assign execute_ctrl1_down_FpuMulPlugin_SUB1_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_SUB1_lane0_1[0];
  assign execute_ctrl1_down_FpuMulPlugin_SUB2_lane0 = _zz_execute_ctrl1_down_FpuMulPlugin_SUB2_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_IS_W_lane0[0];
  assign execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = {(|{_zz_execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0,{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,_zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0}})};
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3;
  assign execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0);
  assign execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0),(|_zz_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1)};
  assign when_ExecuteLanePlugin_l306 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign execute_lane0_ctrls_0_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l306;
  assign when_ExecuteLanePlugin_l306_1 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign execute_lane0_ctrls_1_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l306_1;
  assign when_ExecuteLanePlugin_l306_2 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{((early1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early1_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l306_2 && early1_BranchPlugin_logic_flushPort_payload_self))),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(_zz_when_ExecuteLanePlugin_l306_2_1 && _zz_when_ExecuteLanePlugin_l306_2_2),{_zz_when_ExecuteLanePlugin_l306_2_3,{_zz_when_ExecuteLanePlugin_l306_2_4,_zz_when_ExecuteLanePlugin_l306_2_5}}}}}});
  assign execute_lane0_ctrls_2_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l306_2;
  assign when_ExecuteLanePlugin_l306_3 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}});
  assign execute_lane0_ctrls_3_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l306_3;
  assign when_ExecuteLanePlugin_l306_4 = (|{((late1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late1_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane0) || ((late1_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane0) && late1_BranchPlugin_logic_flushPort_payload_self))),{((late0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late0_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l306_4 && late0_BranchPlugin_logic_flushPort_payload_self))),((LsuPlugin_logic_flushPort_valid && 1'b1) && ((LsuPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l306_4_1 && LsuPlugin_logic_flushPort_payload_self)))}});
  assign execute_lane0_ctrls_4_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l306_4;
  assign execute_lane0_ctrls_5_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_6_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_6_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_7_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_7_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_8_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_8_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_9_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_9_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_10_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_10_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_11_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_11_upIsCancel = 1'b0;
  assign execute_lane0_ctrls_12_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_12_upIsCancel = 1'b0;
  assign execute_lane0_logic_trapPending[0] = (|{((execute_ctrl4_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl4_down_TRAP_lane0),{((execute_ctrl3_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl3_down_TRAP_lane0),{((execute_ctrl2_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl2_down_TRAP_lane0),((execute_ctrl1_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl1_down_TRAP_lane0)}}});
  assign execute_ctrl2_up_COMMIT_lane0 = (! execute_ctrl2_up_TRAP_lane0);
  assign when_FpuFlagsWritebackPlugin_l96 = (! execute_freeze_valid);
  assign WhiteboxerPlugin_logic_csr_access_valid = CsrAccessPlugin_logic_fsm_interface_fire;
  assign WhiteboxerPlugin_logic_csr_access_payload_uopId = CsrAccessPlugin_logic_fsm_interface_uopId;
  assign WhiteboxerPlugin_logic_csr_access_payload_address = _zz_WhiteboxerPlugin_logic_csr_access_payload_address[31 : 20];
  assign WhiteboxerPlugin_logic_csr_access_payload_write = CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  assign WhiteboxerPlugin_logic_csr_access_payload_read = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign WhiteboxerPlugin_logic_csr_access_payload_writeDone = CsrAccessPlugin_logic_fsm_interface_write;
  assign WhiteboxerPlugin_logic_csr_access_payload_readDone = CsrAccessPlugin_logic_fsm_interface_read;
  assign WhiteboxerPlugin_logic_csr_port_valid = WhiteboxerPlugin_logic_csr_access_valid;
  assign WhiteboxerPlugin_logic_csr_port_payload_uopId = WhiteboxerPlugin_logic_csr_access_payload_uopId;
  assign WhiteboxerPlugin_logic_csr_port_payload_address = WhiteboxerPlugin_logic_csr_access_payload_address;
  assign WhiteboxerPlugin_logic_csr_port_payload_write = WhiteboxerPlugin_logic_csr_access_payload_write;
  assign WhiteboxerPlugin_logic_csr_port_payload_read = WhiteboxerPlugin_logic_csr_access_payload_read;
  assign WhiteboxerPlugin_logic_csr_port_payload_writeDone = WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  assign WhiteboxerPlugin_logic_csr_port_payload_readDone = WhiteboxerPlugin_logic_csr_access_payload_readDone;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_valid = lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_valid = lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_valid = lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_valid = lane1_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_payload_uopId = lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_payload_data = lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_valid = lane1_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_payload_uopId = lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_payload_data = lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_valid = lane0_float_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_payload_data = lane0_float_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_6_valid = lane0_float_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_6_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_6_payload_data = lane0_float_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_7_valid = lane0_float_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_7_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_7_payload_data = lane0_float_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_8_valid = lane0_float_WriteBackPlugin_logic_stages_3_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_8_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_3_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_8_payload_data = lane0_float_WriteBackPlugin_logic_stages_3_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_9_valid = lane0_float_WriteBackPlugin_logic_stages_4_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_9_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_4_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_9_payload_data = lane0_float_WriteBackPlugin_logic_stages_4_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_10_valid = lane0_float_WriteBackPlugin_logic_stages_5_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_10_payload_uopId = lane0_float_WriteBackPlugin_logic_stages_5_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_10_payload_data = lane0_float_WriteBackPlugin_logic_stages_5_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_11_valid = FpuPackerPlugin_logic_s2_fpWriter_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_11_payload_uopId = FpuPackerPlugin_logic_s2_fpWriter_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_11_payload_data = FpuPackerPlugin_logic_s2_fpWriter_payload_data;
  assign WhiteboxerPlugin_logic_completions_ports_0_valid = DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_uopId = DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_trap = DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_commit = DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_1_valid = DecoderPlugin_logic_laneLogic_1_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_uopId = DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_trap = DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_commit = DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_2_valid = execute_lane0_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_uopId = execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_trap = execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_commit = execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_3_valid = execute_lane0_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_uopId = execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_trap = execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_commit = execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_4_valid = execute_lane0_logic_completions_onCtrl_2_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_uopId = execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_trap = execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_commit = execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_5_valid = execute_lane0_logic_completions_onCtrl_3_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_uopId = execute_lane0_logic_completions_onCtrl_3_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_trap = execute_lane0_logic_completions_onCtrl_3_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_commit = execute_lane0_logic_completions_onCtrl_3_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_6_valid = execute_lane0_logic_completions_onCtrl_4_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_uopId = execute_lane0_logic_completions_onCtrl_4_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_trap = execute_lane0_logic_completions_onCtrl_4_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_commit = execute_lane0_logic_completions_onCtrl_4_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_7_valid = execute_lane0_logic_completions_onCtrl_5_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_uopId = execute_lane0_logic_completions_onCtrl_5_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_trap = execute_lane0_logic_completions_onCtrl_5_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_commit = execute_lane0_logic_completions_onCtrl_5_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_8_valid = execute_lane0_logic_completions_onCtrl_6_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_8_payload_uopId = execute_lane0_logic_completions_onCtrl_6_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_8_payload_trap = execute_lane0_logic_completions_onCtrl_6_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_8_payload_commit = execute_lane0_logic_completions_onCtrl_6_port_payload_commit;
  assign fetch_logic_flushes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_0_doIt),{_zz_fetch_logic_flushes_0_doIt_1,{_zz_fetch_logic_flushes_0_doIt_2,_zz_fetch_logic_flushes_0_doIt_3}}}}}}}});
  assign fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48 = fetch_logic_flushes_0_doIt;
  assign fetch_logic_flushes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_1_doIt),{_zz_fetch_logic_flushes_1_doIt_1,{_zz_fetch_logic_flushes_1_doIt_2,_zz_fetch_logic_flushes_1_doIt_3}}}}}}}});
  assign fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50 = fetch_logic_flushes_1_doIt;
  always @(*) begin
    execute_lane1_bypasser_integer_RS1_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl2_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[1] = (((execute_ctrl2_up_LANE_SEL_lane1 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl2_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[2] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[3] = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[4] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[5] = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[6] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[7] = (((execute_ctrl5_up_LANE_SEL_lane1 && execute_ctrl5_up_RD_ENABLE_lane1) && (execute_ctrl5_down_RD_PHYS_lane1 == execute_ctrl1_down_RS1_PHYS_lane1)) && (execute_ctrl5_down_RD_RFID_lane1 == execute_ctrl1_down_RS1_RFID_lane1));
    execute_lane1_bypasser_integer_RS1_bypassEnables[8] = 1'b1;
  end

  assign _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 = execute_lane1_bypasser_integer_RS1_bypassEnables;
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[4];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[5];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[6];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[7];
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8 = _zz_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_execute_lane1_bypasser_integer_RS1_sel[0] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane1_bypasser_integer_RS1_sel[1] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1 && (! execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_execute_lane1_bypasser_integer_RS1_sel[2] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2 && (! execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_execute_lane1_bypasser_integer_RS1_sel[3] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3 && (! execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_execute_lane1_bypasser_integer_RS1_sel[4] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 && (! execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3));
    _zz_execute_lane1_bypasser_integer_RS1_sel[5] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5 && (! (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 || execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS1_sel[6] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6 && (! (execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5 || execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS1_sel[7] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7 && (! (execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6 || execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS1_sel[8] = (execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8 && (! (execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7 || execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
  end

  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0});
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4});
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4}});
  assign execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7 = (|{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6,{execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4}}});
  assign execute_lane1_bypasser_integer_RS1_sel = _zz_execute_lane1_bypasser_integer_RS1_sel;
  assign _zz_execute_ctrl1_down_integer_RS1_lane1 = execute_lane1_bypasser_integer_RS1_sel[8 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS1_lane1_1 = ((((_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1 ? execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_1) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_2 ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_3)) | ((_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_4 ? execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_5) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_6 ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_7))) | (((_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_8 ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_9) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_10 ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_11)) | ((_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_12 ? execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_13) | (_zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_14 ? execute_lane1_bypasser_integer_RS1_port_data : _zz__zz_execute_ctrl1_down_integer_RS1_lane1_1_15))));
    if(when_ExecuteLanePlugin_l196_2) begin
      _zz_execute_ctrl1_down_integer_RS1_lane1_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS1_lane1 = _zz_execute_ctrl1_down_integer_RS1_lane1_1;
  assign when_ExecuteLanePlugin_l196_2 = execute_lane1_bypasser_integer_RS1_sel[0];
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit = (execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit && (! (|{execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_1,execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_youngerHits_0})));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit = (execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS1_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit = (execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit && (! (|{execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_1,execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_youngerHits_0})));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits = {execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit,{execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit,execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit}};
  assign _zz_execute_ctrl2_integer_RS1_lane1_bypass = {execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits,(! (|execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits))};
  assign execute_ctrl2_integer_RS1_lane1_bypass = (((_zz_execute_ctrl2_integer_RS1_lane1_bypass[0] ? execute_ctrl2_up_integer_RS1_lane1 : 32'h0) | (_zz_execute_ctrl2_integer_RS1_lane1_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl2_integer_RS1_lane1_bypass[2] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS1_lane1_bypass[3] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0)));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl3_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl3_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit = (execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl3_down_RS1_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl3_down_RS1_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit = (execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits = {execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit,execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit};
  assign _zz_execute_ctrl3_integer_RS1_lane1_bypass = {execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits,(! (|execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits))};
  assign execute_ctrl3_integer_RS1_lane1_bypass = (((_zz_execute_ctrl3_integer_RS1_lane1_bypass[0] ? execute_ctrl3_up_integer_RS1_lane1 : 32'h0) | (_zz_execute_ctrl3_integer_RS1_lane1_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_execute_ctrl3_integer_RS1_lane1_bypass[2] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane1_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign execute_lane1_bypasser_integer_RS2_port_address = execute_ctrl0_down_RS2_PHYS_lane1[4 : 0];
  always @(*) begin
    execute_lane1_bypasser_integer_RS2_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl2_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[1] = (((execute_ctrl2_up_LANE_SEL_lane1 && execute_ctrl2_up_RD_ENABLE_lane1) && (execute_ctrl2_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl2_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[2] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[3] = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[4] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[5] = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[6] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl5_down_RD_RFID_lane0 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[7] = (((execute_ctrl5_up_LANE_SEL_lane1 && execute_ctrl5_up_RD_ENABLE_lane1) && (execute_ctrl5_down_RD_PHYS_lane1 == execute_ctrl1_down_RS2_PHYS_lane1)) && (execute_ctrl5_down_RD_RFID_lane1 == execute_ctrl1_down_RS2_RFID_lane1));
    execute_lane1_bypasser_integer_RS2_bypassEnables[8] = 1'b1;
  end

  assign _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 = execute_lane1_bypasser_integer_RS2_bypassEnables;
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[4];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[5];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[6];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[7];
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8 = _zz_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_execute_lane1_bypasser_integer_RS2_sel[0] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane1_bypasser_integer_RS2_sel[1] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1 && (! execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_execute_lane1_bypasser_integer_RS2_sel[2] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2 && (! execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_execute_lane1_bypasser_integer_RS2_sel[3] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3 && (! execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_execute_lane1_bypasser_integer_RS2_sel[4] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 && (! execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3));
    _zz_execute_lane1_bypasser_integer_RS2_sel[5] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5 && (! (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 || execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS2_sel[6] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6 && (! (execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5 || execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS2_sel[7] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7 && (! (execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6 || execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_execute_lane1_bypasser_integer_RS2_sel[8] = (execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8 && (! (execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7 || execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
  end

  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0});
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4});
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4}});
  assign execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7 = (|{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6,{execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4}}});
  assign execute_lane1_bypasser_integer_RS2_sel = _zz_execute_lane1_bypasser_integer_RS2_sel;
  assign _zz_execute_ctrl1_down_integer_RS2_lane1 = execute_lane1_bypasser_integer_RS2_sel[8 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS2_lane1_1 = ((((_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1 ? execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_1) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_2 ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_3)) | ((_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_4 ? execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_5) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_6 ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_7))) | (((_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_8 ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_9) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_10 ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_11)) | ((_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_12 ? execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_13) | (_zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_14 ? execute_lane1_bypasser_integer_RS2_port_data : _zz__zz_execute_ctrl1_down_integer_RS2_lane1_1_15))));
    if(when_ExecuteLanePlugin_l196_3) begin
      _zz_execute_ctrl1_down_integer_RS2_lane1_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS2_lane1 = _zz_execute_ctrl1_down_integer_RS2_lane1_1;
  assign when_ExecuteLanePlugin_l196_3 = execute_lane1_bypasser_integer_RS2_sel[0];
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit = (execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit && (! (|{execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_1,execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_youngerHits_0})));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit = (execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0 = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane0 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1 = (((execute_ctrl3_up_LANE_SEL_lane1 && execute_ctrl3_up_RD_ENABLE_lane1) && (execute_ctrl3_down_RD_PHYS_lane1 == execute_ctrl2_down_RS2_PHYS_lane1)) && (execute_ctrl3_down_RD_RFID_lane1 == execute_ctrl2_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit = (execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit && (! (|{execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_1,execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_youngerHits_0})));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits = {execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit,{execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit,execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit}};
  assign _zz_execute_ctrl2_integer_RS2_lane1_bypass = {execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits,(! (|execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits))};
  assign execute_ctrl2_integer_RS2_lane1_bypass = (((_zz_execute_ctrl2_integer_RS2_lane1_bypass[0] ? execute_ctrl2_up_integer_RS2_lane1 : 32'h0) | (_zz_execute_ctrl2_integer_RS2_lane1_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl2_integer_RS2_lane1_bypass[2] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl2_integer_RS2_lane1_bypass[3] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0)));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl3_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane0 == execute_ctrl3_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit = (execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit = (((execute_ctrl4_up_LANE_SEL_lane1 && execute_ctrl4_up_RD_ENABLE_lane1) && (execute_ctrl4_down_RD_PHYS_lane1 == execute_ctrl3_down_RS2_PHYS_lane1)) && (execute_ctrl4_down_RD_RFID_lane1 == execute_ctrl3_down_RS2_RFID_lane1));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit = (execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits = {execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit,execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit};
  assign _zz_execute_ctrl3_integer_RS2_lane1_bypass = {execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits,(! (|execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits))};
  assign execute_ctrl3_integer_RS2_lane1_bypass = (((_zz_execute_ctrl3_integer_RS2_lane1_bypass[0] ? execute_ctrl3_up_integer_RS2_lane1 : 32'h0) | (_zz_execute_ctrl3_integer_RS2_lane1_bypass[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_execute_ctrl3_integer_RS2_lane1_bypass[2] ? execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane1_logic_completions_onCtrl_0_port_valid = (((execute_ctrl2_down_LANE_SEL_lane1 && execute_ctrl2_down_isReady) && (! execute_lane1_ctrls_2_downIsCancel)) && execute_ctrl2_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1);
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_trap = execute_ctrl2_down_TRAP_lane1;
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_commit = execute_ctrl2_down_COMMIT_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_valid = (((execute_ctrl4_down_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_downIsCancel)) && execute_ctrl4_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1);
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_trap = execute_ctrl4_down_TRAP_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_commit = execute_ctrl4_down_COMMIT_lane1;
  assign execute_lane1_logic_decoding_decodingBits = {execute_ctrl1_down_lane1_LAYER_SEL_lane1,execute_ctrl1_down_Decode_UOP_lane1};
  always @(*) begin
    execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = _zz_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = _zz_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000010) == 33'h0);
  always @(*) begin
    execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = _zz_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000000004) == 33'h000000004);
  always @(*) begin
    execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = _zz_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000000) == 33'h100000000);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_2_lane1 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_COMPLETION_AT_2_lane1 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000000) == 33'h0);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_4_lane1 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_COMPLETION_AT_4_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = _zz_execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1[0];
    if(execute_ctrl1_down_TRAP_lane1) begin
      execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000006000) == 33'h0);
  assign execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000006004) == 33'h000002000);
  assign execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000003000) == 33'h000002000);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000004000) == 33'h0);
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000001000) == 33'h000001000);
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1 = {(|{_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1,{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1}}),(|{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1,_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1}})};
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  assign _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  assign execute_ctrl1_down_SrcStageables_REVERT_lane1 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane1[0];
  assign execute_ctrl1_down_SrcStageables_ZERO_lane1 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane1[0];
  assign execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h000000044) == 33'h000000004));
  assign _zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000000024) == 33'h0);
  assign execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1 = {(|_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1),(|_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1)};
  assign execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1 = _zz_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1[0];
  assign execute_ctrl1_down_BYPASSED_AT_2_lane1 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane1[0];
  assign execute_ctrl1_down_BYPASSED_AT_3_lane1 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane1_1[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1[0];
  assign execute_ctrl1_down_SrcStageables_UNSIGNED_lane1 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1[0];
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1 = {(|((execute_lane1_logic_decoding_decodingBits & 33'h00000000c) == 33'h000000004)),(|((execute_lane1_logic_decoding_decodingBits & 33'h000000008) == 33'h000000008))};
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1;
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  assign execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2;
  assign execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1[0];
  assign execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1[0];
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3 = {(|{_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1,{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1}}),(|{_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1,_zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1}})};
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3;
  assign _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  assign execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4;
  assign execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = (|_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1);
  assign execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = {(|_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1),(|_zz_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1)};
  assign when_ExecuteLanePlugin_l306_5 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign execute_lane1_ctrls_0_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l306_5;
  assign when_ExecuteLanePlugin_l306_6 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign execute_lane1_ctrls_1_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l306_6;
  assign when_ExecuteLanePlugin_l306_7 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{((early1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early1_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl2_down_LANE_AGE_lane1) || ((early1_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl2_down_LANE_AGE_lane1) && early1_BranchPlugin_logic_flushPort_payload_self))),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{((early0_EnvPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l306_7) && (_zz_when_ExecuteLanePlugin_l306_7_1 || _zz_when_ExecuteLanePlugin_l306_7_2)),{(_zz_when_ExecuteLanePlugin_l306_7_3 && _zz_when_ExecuteLanePlugin_l306_7_4),{_zz_when_ExecuteLanePlugin_l306_7_5,_zz_when_ExecuteLanePlugin_l306_7_6}}}}}});
  assign execute_lane1_ctrls_2_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l306_7;
  assign when_ExecuteLanePlugin_l306_8 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}});
  assign execute_lane1_ctrls_3_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l306_8;
  assign when_ExecuteLanePlugin_l306_9 = (|{((late1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late1_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane1) || ((late1_BranchPlugin_logic_flushPort_payload_laneAge == execute_ctrl4_down_LANE_AGE_lane1) && late1_BranchPlugin_logic_flushPort_payload_self))),{((late0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late0_BranchPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane1) || (_zz_when_ExecuteLanePlugin_l306_9 && late0_BranchPlugin_logic_flushPort_payload_self))),((LsuPlugin_logic_flushPort_valid && 1'b1) && ((LsuPlugin_logic_flushPort_payload_laneAge < execute_ctrl4_down_LANE_AGE_lane1) || (_zz_when_ExecuteLanePlugin_l306_9_1 && LsuPlugin_logic_flushPort_payload_self)))}});
  assign execute_lane1_ctrls_4_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l306_9;
  assign execute_lane1_ctrls_5_downIsCancel = 1'b0;
  assign execute_lane1_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane1_logic_trapPending[0] = (|{((execute_ctrl4_up_LANE_SEL_lane1 && 1'b1) && execute_ctrl4_down_TRAP_lane1),{((execute_ctrl3_up_LANE_SEL_lane1 && 1'b1) && execute_ctrl3_down_TRAP_lane1),{((execute_ctrl2_up_LANE_SEL_lane1 && 1'b1) && execute_ctrl2_down_TRAP_lane1),((execute_ctrl1_up_LANE_SEL_lane1 && 1'b1) && execute_ctrl1_down_TRAP_lane1)}}});
  assign execute_ctrl2_up_COMMIT_lane1 = (! execute_ctrl2_up_TRAP_lane1);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (|lane0_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = lane0_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = lane0_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_uopId = lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_valid = (|lane1_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_address = lane1_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_data = lane1_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_uopId = lane1_integer_WriteBackPlugin_logic_write_port_uopId;
  assign execute_lane1_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  assign execute_lane0_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  assign execute_lane0_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  assign execute_lane1_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_initalizer_counter[4:0];
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
    if(when_RegFilePlugin_l132) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = 32'h0;
    end
  end

  assign integer_RegFilePlugin_logic_initalizer_done = integer_RegFilePlugin_logic_initalizer_counter[5];
  assign when_RegFilePlugin_l132 = (! integer_RegFilePlugin_logic_initalizer_done);
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_uopId = integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  assign integer_write_1_valid = integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  assign integer_write_1_address = integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  assign integer_write_1_data = integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  assign integer_write_1_uopId = integer_RegFilePlugin_logic_writeMerges_1_bus_uopId;
  assign float_RegFilePlugin_logic_writeMerges_0_bus_valid = (|lane0_float_WriteBackPlugin_logic_write_port_valid);
  assign float_RegFilePlugin_logic_writeMerges_0_bus_address = lane0_float_WriteBackPlugin_logic_write_port_address;
  assign float_RegFilePlugin_logic_writeMerges_0_bus_data = lane0_float_WriteBackPlugin_logic_write_port_data;
  assign float_RegFilePlugin_logic_writeMerges_0_bus_uopId = lane0_float_WriteBackPlugin_logic_write_port_uopId;
  assign execute_lane0_bypasser_float_RS1_port_data = float_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  assign execute_lane0_bypasser_float_RS2_port_data = float_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  assign execute_lane0_bypasser_float_RS3_port_data = float_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  always @(*) begin
    float_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = float_RegFilePlugin_logic_writeMerges_0_bus_valid;
    if(when_RegFilePlugin_l132_1) begin
      float_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    float_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = float_RegFilePlugin_logic_writeMerges_0_bus_address;
    if(when_RegFilePlugin_l132_1) begin
      float_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = float_RegFilePlugin_logic_initalizer_counter[4:0];
    end
  end

  always @(*) begin
    float_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = float_RegFilePlugin_logic_writeMerges_0_bus_data;
    if(when_RegFilePlugin_l132_1) begin
      float_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = 64'h0;
    end
  end

  assign float_RegFilePlugin_logic_initalizer_done = float_RegFilePlugin_logic_initalizer_counter[5];
  assign when_RegFilePlugin_l132_1 = (! float_RegFilePlugin_logic_initalizer_done);
  assign float_write_0_valid = float_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign float_write_0_address = float_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign float_write_0_data = float_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign float_write_0_uopId = float_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  assign execute_freeze_valid = (|{CsrAccessPlugin_logic_fsm_inject_freeze,{FpuSqrtPlugin_logic_onExecute_freeze,{FpuF2iPlugin_logic_onResult_halfRater_freezeIt,{FpuUnpackerPlugin_logic_onCvt_freezeIt,{FpuUnpack_RS3_normalizer_freezeIt,{FpuUnpack_RS2_normalizer_freezeIt,{FpuUnpack_RS1_normalizer_freezeIt,{FpuPackerPlugin_logic_s1_subnormal_freezeIt,{LsuPlugin_logic_onCtrl_rva_freezeIt,{LsuPlugin_logic_onCtrl_io_freezeIt,early0_DivPlugin_logic_processing_freeze}}}}}}}}}});
  assign execute_ctrl12_down_ready = (! execute_freeze_valid);
  assign WhiteboxerPlugin_logic_completions_ports_9_valid = execute_lane1_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_9_payload_uopId = execute_lane1_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_9_payload_trap = execute_lane1_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_9_payload_commit = execute_lane1_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_10_valid = execute_lane1_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_10_payload_uopId = execute_lane1_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_10_payload_trap = execute_lane1_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_10_payload_commit = execute_lane1_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_0 = ((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane0) && (execute_ctrl4_down_LANE_AGE_lane0 == 1'b0));
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_1 = ((((execute_ctrl4_down_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane1) && (execute_ctrl4_down_LANE_AGE_lane1 == 1'b0));
  assign WhiteboxerPlugin_logic_commits_ports_0_valid = (|{WhiteboxerPlugin_logic_commits_ports_0_oh_1,WhiteboxerPlugin_logic_commits_ports_0_oh_0});
  assign WhiteboxerPlugin_logic_commits_ports_0_pc = ((WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_PC_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_0_oh_1 ? execute_ctrl4_down_PC_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_0_uop = ((WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_Decode_UOP_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_0_oh_1 ? execute_ctrl4_down_Decode_UOP_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_1_oh_0 = ((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane0) && (execute_ctrl4_down_LANE_AGE_lane0 == 1'b1));
  assign WhiteboxerPlugin_logic_commits_ports_1_oh_1 = ((((execute_ctrl4_down_LANE_SEL_lane1 && execute_ctrl4_down_isReady) && (! execute_lane1_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane1) && (execute_ctrl4_down_LANE_AGE_lane1 == 1'b1));
  assign WhiteboxerPlugin_logic_commits_ports_1_valid = (|{WhiteboxerPlugin_logic_commits_ports_1_oh_1,WhiteboxerPlugin_logic_commits_ports_1_oh_0});
  assign WhiteboxerPlugin_logic_commits_ports_1_pc = ((WhiteboxerPlugin_logic_commits_ports_1_oh_0 ? execute_ctrl4_down_PC_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_1_oh_1 ? execute_ctrl4_down_PC_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_1_uop = ((WhiteboxerPlugin_logic_commits_ports_1_oh_0 ? execute_ctrl4_down_Decode_UOP_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_1_oh_1 ? execute_ctrl4_down_Decode_UOP_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_valid = BtbPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self = BtbPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_valid = LsuPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId = LsuPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_laneAge = LsuPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self = LsuPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_valid = early0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId = early0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_laneAge = early0_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self = early0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_valid = CsrAccessPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId = CsrAccessPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_laneAge = CsrAccessPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self = CsrAccessPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_valid = early0_EnvPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId = early0_EnvPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_laneAge = early0_EnvPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self = early0_EnvPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_valid = late0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId = late0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_laneAge = late0_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self = late0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_valid = early1_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_uopId = early1_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_laneAge = early1_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_self = early1_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_valid = late1_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_uopId = late1_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_laneAge = late1_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_self = late1_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_valid = DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_uopId = DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_laneAge = DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_self = DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_valid = DecoderPlugin_logic_laneLogic_1_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_uopId = DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_laneAge = DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_self = DecoderPlugin_logic_laneLogic_1_flushPort_payload_self;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid = late0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice = late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget = late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken = late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch = late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush = late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop = late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget = late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history = late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId = late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign WhiteboxerPlugin_logic_prediction_learns_0_valid = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_taken = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_history = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_valid = late1_BranchPlugin_logic_jumpLogic_learn_valid;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice = late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget = late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken = late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch = late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush = late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop = late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget = late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history = late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId = late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign WhiteboxerPlugin_logic_prediction_learns_1_valid = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_pcOnLastSlice = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_pcTarget = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_taken = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isBranch = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isPush = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isPop = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_badPredictedTarget = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_history = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_uopId = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late1_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign WhiteboxerPlugin_logic_loadExecute_fire = (((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_AguPlugin_LOAD_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0)) && (! execute_ctrl4_down_TRAP_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign WhiteboxerPlugin_logic_loadExecute_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  always @(*) begin
    WhiteboxerPlugin_logic_loadExecute_data = {32'd0, lane0_IntFormatPlugin_logic_stages_1_wb_payload};
    if(LsuPlugin_logic_fpwb_valid) begin
      WhiteboxerPlugin_logic_loadExecute_data = _zz_WhiteboxerPlugin_logic_loadExecute_data;
    end
  end

  assign WhiteboxerPlugin_logic_storeCommit_fire = LsuPlugin_logic_onWb_storeFire;
  assign WhiteboxerPlugin_logic_storeCommit_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_address = execute_ctrl4_down_MMU_TRANSLATED_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_amo = 1'b0;
  assign WhiteboxerPlugin_logic_storeConditional_fire = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && (execute_ctrl4_down_AguPlugin_ATOMIC_lane0 && (! execute_ctrl4_down_AguPlugin_LOAD_lane0))) && (! execute_ctrl4_down_TRAP_lane0));
  assign WhiteboxerPlugin_logic_storeConditional_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeConditional_miss = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  assign WhiteboxerPlugin_logic_storeBroadcast_fire = LsuPlugin_logic_onWb_storeBroadcast;
  assign WhiteboxerPlugin_logic_storeBroadcast_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign TrapPlugin_logic_initHold = (|{(! float_RegFilePlugin_logic_initalizer_done),{(! CsrRamPlugin_logic_flush_done),{1'b0,{((! LsuL1Plugin_logic_initializer_done) || 1'b0),{(! integer_RegFilePlugin_logic_initalizer_done),{(FetchL1Plugin_logic_invalidate_firstEver || _zz_TrapPlugin_logic_initHold),{_zz_TrapPlugin_logic_initHold_1,_zz_TrapPlugin_logic_initHold_2}}}}}}});
  assign WhiteboxerPlugin_logic_wfi = TrapPlugin_logic_harts_0_trap_fsm_wfi;
  assign WhiteboxerPlugin_logic_perf_executeFreezed = execute_freeze_valid;
  assign WhiteboxerPlugin_logic_perf_dispatchHazards = (|{(DispatchPlugin_logic_candidates_2_ctx_valid && (! DispatchPlugin_logic_candidates_2_fire)),{(DispatchPlugin_logic_candidates_1_ctx_valid && (! DispatchPlugin_logic_candidates_1_fire)),(DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_fire))}});
  assign WhiteboxerPlugin_logic_perf_candidatesCount = _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  assign WhiteboxerPlugin_logic_perf_dispatchFeedCount = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_executeFreezed) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_executeFreezedCounter = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_dispatchHazards) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  assign when_Utils_l593 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b00);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b0;
    if(when_Utils_l593) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  assign when_Utils_l593_1 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b01);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b0;
    if(when_Utils_l593_1) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  assign when_Utils_l593_2 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b10);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = 1'b0;
    if(when_Utils_l593_2) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2;
  assign when_Utils_l593_3 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b11);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = 1'b0;
    if(when_Utils_l593_3) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2;
  assign when_Utils_l593_4 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b00);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b0;
    if(when_Utils_l593_4) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  assign when_Utils_l593_5 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b01);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b0;
    if(when_Utils_l593_5) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  assign when_Utils_l593_6 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b10);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = 1'b0;
    if(when_Utils_l593_6) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2;
  assign WhiteboxerPlugin_logic_trap_ports_0_valid = TrapPlugin_logic_harts_0_trap_whitebox_trap;
  assign WhiteboxerPlugin_logic_trap_ports_0_interrupt = TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  assign WhiteboxerPlugin_logic_trap_ports_0_cause = TrapPlugin_logic_harts_0_trap_whitebox_code;
  assign fetch_logic_ctrls_2_up_forgetOne = (|fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50);
  assign fetch_logic_ctrls_2_up_cancel = (|fetch_logic_flushes_1_doIt);
  assign fetch_logic_ctrls_1_up_forgetOne = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_up_cancel = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_0_down_ready = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_down_ready = fetch_logic_ctrls_2_up_ready;
  always @(*) begin
    fetch_logic_ctrls_0_down_valid = fetch_logic_ctrls_0_up_valid;
    if(when_CtrlLink_l191) begin
      fetch_logic_ctrls_0_down_valid = 1'b0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_0_up_ready = fetch_logic_ctrls_0_down_isReady;
    if(when_CtrlLink_l191) begin
      fetch_logic_ctrls_0_up_ready = 1'b0;
    end
  end

  assign when_CtrlLink_l191 = (|{fetch_logic_ctrls_0_haltRequest_PcPlugin_l133,{fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200,{fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297,fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217}}});
  assign fetch_logic_ctrls_0_down_Fetch_WORD_PC = fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_0_down_Fetch_PC_FAULT = fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_0_down_Fetch_ID = fetch_logic_ctrls_0_up_Fetch_ID;
  always @(*) begin
    fetch_logic_ctrls_1_down_valid = fetch_logic_ctrls_1_up_valid;
    if(when_CtrlLink_l198) begin
      fetch_logic_ctrls_1_down_valid = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_up_ready = fetch_logic_ctrls_1_down_isReady;
  assign when_CtrlLink_l198 = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_down_Fetch_WORD_PC = fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_1_down_Fetch_PC_FAULT = fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_1_down_Fetch_ID = fetch_logic_ctrls_1_up_Fetch_ID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  assign fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS = fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  assign fetch_logic_ctrls_2_down_valid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_ready = fetch_logic_ctrls_2_down_isReady;
  assign fetch_logic_ctrls_2_down_Fetch_WORD_PC = fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_2_down_Fetch_PC_FAULT = fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_2_down_Fetch_ID = fetch_logic_ctrls_2_up_Fetch_ID;
  assign fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  assign fetch_logic_ctrls_2_down_MMU_TRANSLATED = fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED = fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE = fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC = fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  assign fetch_logic_ctrls_2_down_MMU_REFILL = fetch_logic_ctrls_2_up_MMU_REFILL;
  assign fetch_logic_ctrls_2_down_MMU_HAZARD = fetch_logic_ctrls_2_up_MMU_HAZARD;
  assign fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE = fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  assign fetch_logic_ctrls_2_down_MMU_PAGE_FAULT = fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  assign fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT = fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  assign fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION = fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  always @(*) begin
    decode_ctrls_0_down_ready = decode_ctrls_1_up_ready;
    if(when_StageLink_l71_3) begin
      decode_ctrls_0_down_ready = 1'b1;
    end
  end

  assign when_StageLink_l71_3 = (! decode_ctrls_1_up_isValid);
  assign when_DecodePipelinePlugin_l70 = ((! decode_ctrls_1_up_isReady) && decode_ctrls_1_lane0_upIsCancel);
  assign when_DecodePipelinePlugin_l70_1 = ((! decode_ctrls_1_up_isReady) && decode_ctrls_1_lane1_upIsCancel);
  assign decode_ctrls_0_down_valid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_ready = decode_ctrls_0_down_isReady;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_0 = decode_ctrls_0_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0 = decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign decode_ctrls_0_down_PC_0 = decode_ctrls_0_up_PC_0;
  assign decode_ctrls_0_down_Decode_DOP_ID_0 = decode_ctrls_0_up_Decode_DOP_ID_0;
  assign decode_ctrls_0_down_Fetch_ID_0 = decode_ctrls_0_up_Fetch_ID_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3;
  assign decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_0_down_TRAP_0 = decode_ctrls_0_up_TRAP_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_0_down_Prediction_ALIGN_REDO_0 = decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_1 = decode_ctrls_0_up_Decode_INSTRUCTION_1;
  assign decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1 = decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1 = decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1 = decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign decode_ctrls_0_down_PC_1 = decode_ctrls_0_up_PC_1;
  assign decode_ctrls_0_down_Decode_DOP_ID_1 = decode_ctrls_0_up_Decode_DOP_ID_1;
  assign decode_ctrls_0_down_Fetch_ID_1 = decode_ctrls_0_up_Fetch_ID_1;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3;
  assign decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1 = decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1;
  assign decode_ctrls_0_down_TRAP_1 = decode_ctrls_0_up_TRAP_1;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign decode_ctrls_0_down_Prediction_ALIGN_REDO_1 = decode_ctrls_0_up_Prediction_ALIGN_REDO_1;
  assign decode_ctrls_1_down_valid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_ready = decode_ctrls_1_down_isReady;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_0 = decode_ctrls_1_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0 = decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign decode_ctrls_1_down_PC_0 = decode_ctrls_1_up_PC_0;
  assign decode_ctrls_1_down_Decode_DOP_ID_0 = decode_ctrls_1_up_Decode_DOP_ID_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3;
  assign decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_1_down_Prediction_ALIGN_REDO_0 = decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_1 = decode_ctrls_1_up_Decode_INSTRUCTION_1;
  assign decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1 = decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1 = decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1 = decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign decode_ctrls_1_down_PC_1 = decode_ctrls_1_up_PC_1;
  assign decode_ctrls_1_down_Decode_DOP_ID_1 = decode_ctrls_1_up_Decode_DOP_ID_1;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3;
  assign decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1 = decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign decode_ctrls_1_down_Prediction_ALIGN_REDO_1 = decode_ctrls_1_up_Prediction_ALIGN_REDO_1;
  assign execute_ctrl0_down_ready = execute_ctrl1_up_ready;
  assign execute_ctrl1_down_ready = execute_ctrl2_up_ready;
  assign execute_ctrl2_down_ready = execute_ctrl3_up_ready;
  assign execute_ctrl3_down_ready = execute_ctrl4_up_ready;
  assign execute_ctrl4_down_ready = execute_ctrl5_up_ready;
  assign execute_ctrl5_down_ready = execute_ctrl6_up_ready;
  assign execute_ctrl6_down_ready = execute_ctrl7_up_ready;
  assign execute_ctrl7_down_ready = execute_ctrl8_up_ready;
  assign execute_ctrl8_down_ready = execute_ctrl9_up_ready;
  assign execute_ctrl9_down_ready = execute_ctrl10_up_ready;
  assign execute_ctrl10_down_ready = execute_ctrl11_up_ready;
  assign execute_ctrl11_down_ready = execute_ctrl12_up_ready;
  assign execute_ctrl0_up_ready = execute_ctrl0_down_isReady;
  assign execute_ctrl0_down_Decode_UOP_lane0 = execute_ctrl0_up_Decode_UOP_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  assign execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl0_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl0_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0 = execute_ctrl0_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  assign execute_ctrl0_down_PC_lane0 = execute_ctrl0_up_PC_lane0;
  assign execute_ctrl0_down_TRAP_lane0 = execute_ctrl0_up_TRAP_lane0;
  assign execute_ctrl0_down_Decode_UOP_ID_lane0 = execute_ctrl0_up_Decode_UOP_ID_lane0;
  assign execute_ctrl0_down_RS1_ENABLE_lane0 = execute_ctrl0_up_RS1_ENABLE_lane0;
  assign execute_ctrl0_down_RS1_RFID_lane0 = execute_ctrl0_up_RS1_RFID_lane0;
  assign execute_ctrl0_down_RS1_PHYS_lane0 = execute_ctrl0_up_RS1_PHYS_lane0;
  assign execute_ctrl0_down_RS2_ENABLE_lane0 = execute_ctrl0_up_RS2_ENABLE_lane0;
  assign execute_ctrl0_down_RS2_RFID_lane0 = execute_ctrl0_up_RS2_RFID_lane0;
  assign execute_ctrl0_down_RS2_PHYS_lane0 = execute_ctrl0_up_RS2_PHYS_lane0;
  assign execute_ctrl0_down_RD_RFID_lane0 = execute_ctrl0_up_RD_RFID_lane0;
  assign execute_ctrl0_down_RD_PHYS_lane0 = execute_ctrl0_up_RD_PHYS_lane0;
  assign execute_ctrl0_down_RS3_ENABLE_lane0 = execute_ctrl0_up_RS3_ENABLE_lane0;
  assign execute_ctrl0_down_RS3_RFID_lane0 = execute_ctrl0_up_RS3_RFID_lane0;
  assign execute_ctrl0_down_RS3_PHYS_lane0 = execute_ctrl0_up_RS3_PHYS_lane0;
  assign execute_ctrl0_down_LANE_AGE_lane0 = execute_ctrl0_up_LANE_AGE_lane0;
  assign execute_ctrl0_down_COMPLETED_lane0 = execute_ctrl0_up_COMPLETED_lane0;
  assign execute_ctrl0_down_lane0_LAYER_SEL_lane0 = execute_ctrl0_up_lane0_LAYER_SEL_lane0;
  assign execute_ctrl0_down_Decode_UOP_lane1 = execute_ctrl0_up_Decode_UOP_lane1;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1 = execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1;
  assign execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign execute_ctrl0_down_PC_lane1 = execute_ctrl0_up_PC_lane1;
  assign execute_ctrl0_down_TRAP_lane1 = execute_ctrl0_up_TRAP_lane1;
  assign execute_ctrl0_down_Decode_UOP_ID_lane1 = execute_ctrl0_up_Decode_UOP_ID_lane1;
  assign execute_ctrl0_down_RS1_RFID_lane1 = execute_ctrl0_up_RS1_RFID_lane1;
  assign execute_ctrl0_down_RS1_PHYS_lane1 = execute_ctrl0_up_RS1_PHYS_lane1;
  assign execute_ctrl0_down_RS2_RFID_lane1 = execute_ctrl0_up_RS2_RFID_lane1;
  assign execute_ctrl0_down_RS2_PHYS_lane1 = execute_ctrl0_up_RS2_PHYS_lane1;
  assign execute_ctrl0_down_RD_RFID_lane1 = execute_ctrl0_up_RD_RFID_lane1;
  assign execute_ctrl0_down_RD_PHYS_lane1 = execute_ctrl0_up_RD_PHYS_lane1;
  assign execute_ctrl0_down_LANE_AGE_lane1 = execute_ctrl0_up_LANE_AGE_lane1;
  assign execute_ctrl0_down_COMPLETED_lane1 = execute_ctrl0_up_COMPLETED_lane1;
  assign execute_ctrl0_down_lane1_LAYER_SEL_lane1 = execute_ctrl0_up_lane1_LAYER_SEL_lane1;
  assign execute_ctrl1_up_ready = execute_ctrl1_down_isReady;
  assign execute_ctrl1_down_Decode_UOP_lane0 = execute_ctrl1_up_Decode_UOP_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  assign execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl1_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0 = execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
  assign execute_ctrl1_down_PC_lane0 = execute_ctrl1_up_PC_lane0;
  assign execute_ctrl1_down_TRAP_lane0 = execute_ctrl1_up_TRAP_lane0;
  assign execute_ctrl1_down_Decode_UOP_ID_lane0 = execute_ctrl1_up_Decode_UOP_ID_lane0;
  assign execute_ctrl1_down_RS1_ENABLE_lane0 = execute_ctrl1_up_RS1_ENABLE_lane0;
  assign execute_ctrl1_down_RS1_RFID_lane0 = execute_ctrl1_up_RS1_RFID_lane0;
  assign execute_ctrl1_down_RS1_PHYS_lane0 = execute_ctrl1_up_RS1_PHYS_lane0;
  assign execute_ctrl1_down_RS2_ENABLE_lane0 = execute_ctrl1_up_RS2_ENABLE_lane0;
  assign execute_ctrl1_down_RS2_RFID_lane0 = execute_ctrl1_up_RS2_RFID_lane0;
  assign execute_ctrl1_down_RS2_PHYS_lane0 = execute_ctrl1_up_RS2_PHYS_lane0;
  assign execute_ctrl1_down_RD_RFID_lane0 = execute_ctrl1_up_RD_RFID_lane0;
  assign execute_ctrl1_down_RD_PHYS_lane0 = execute_ctrl1_up_RD_PHYS_lane0;
  assign execute_ctrl1_down_RS3_ENABLE_lane0 = execute_ctrl1_up_RS3_ENABLE_lane0;
  assign execute_ctrl1_down_RS3_RFID_lane0 = execute_ctrl1_up_RS3_RFID_lane0;
  assign execute_ctrl1_down_RS3_PHYS_lane0 = execute_ctrl1_up_RS3_PHYS_lane0;
  assign execute_ctrl1_down_LANE_AGE_lane0 = execute_ctrl1_up_LANE_AGE_lane0;
  assign execute_ctrl1_down_COMPLETED_lane0 = execute_ctrl1_up_COMPLETED_lane0;
  assign execute_ctrl1_down_lane0_LAYER_SEL_lane0 = execute_ctrl1_up_lane0_LAYER_SEL_lane0;
  assign execute_ctrl1_down_Decode_UOP_lane1 = execute_ctrl1_up_Decode_UOP_lane1;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1 = execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1;
  assign execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign execute_ctrl1_down_PC_lane1 = execute_ctrl1_up_PC_lane1;
  assign execute_ctrl1_down_TRAP_lane1 = execute_ctrl1_up_TRAP_lane1;
  assign execute_ctrl1_down_Decode_UOP_ID_lane1 = execute_ctrl1_up_Decode_UOP_ID_lane1;
  assign execute_ctrl1_down_RS1_RFID_lane1 = execute_ctrl1_up_RS1_RFID_lane1;
  assign execute_ctrl1_down_RS1_PHYS_lane1 = execute_ctrl1_up_RS1_PHYS_lane1;
  assign execute_ctrl1_down_RS2_RFID_lane1 = execute_ctrl1_up_RS2_RFID_lane1;
  assign execute_ctrl1_down_RS2_PHYS_lane1 = execute_ctrl1_up_RS2_PHYS_lane1;
  assign execute_ctrl1_down_RD_RFID_lane1 = execute_ctrl1_up_RD_RFID_lane1;
  assign execute_ctrl1_down_RD_PHYS_lane1 = execute_ctrl1_up_RD_PHYS_lane1;
  assign execute_ctrl1_down_LANE_AGE_lane1 = execute_ctrl1_up_LANE_AGE_lane1;
  assign execute_ctrl1_down_COMPLETED_lane1 = execute_ctrl1_up_COMPLETED_lane1;
  assign execute_ctrl1_down_lane1_LAYER_SEL_lane1 = execute_ctrl1_up_lane1_LAYER_SEL_lane1;
  assign execute_ctrl1_down_AguPlugin_SIZE_lane0 = execute_ctrl1_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_up_ready = execute_ctrl2_down_isReady;
  assign execute_ctrl2_down_Decode_UOP_lane0 = execute_ctrl2_up_Decode_UOP_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  assign execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl2_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl2_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl2_down_PC_lane0 = execute_ctrl2_up_PC_lane0;
  assign execute_ctrl2_down_Decode_UOP_ID_lane0 = execute_ctrl2_up_Decode_UOP_ID_lane0;
  assign execute_ctrl2_down_RS1_RFID_lane0 = execute_ctrl2_up_RS1_RFID_lane0;
  assign execute_ctrl2_down_RS1_PHYS_lane0 = execute_ctrl2_up_RS1_PHYS_lane0;
  assign execute_ctrl2_down_RS2_RFID_lane0 = execute_ctrl2_up_RS2_RFID_lane0;
  assign execute_ctrl2_down_RS2_PHYS_lane0 = execute_ctrl2_up_RS2_PHYS_lane0;
  assign execute_ctrl2_down_RD_RFID_lane0 = execute_ctrl2_up_RD_RFID_lane0;
  assign execute_ctrl2_down_RD_PHYS_lane0 = execute_ctrl2_up_RD_PHYS_lane0;
  assign execute_ctrl2_down_RS3_RFID_lane0 = execute_ctrl2_up_RS3_RFID_lane0;
  assign execute_ctrl2_down_LANE_AGE_lane0 = execute_ctrl2_up_LANE_AGE_lane0;
  assign execute_ctrl2_down_Decode_UOP_lane1 = execute_ctrl2_up_Decode_UOP_lane1;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1 = execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1;
  assign execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign execute_ctrl2_down_PC_lane1 = execute_ctrl2_up_PC_lane1;
  assign execute_ctrl2_down_TRAP_lane1 = execute_ctrl2_up_TRAP_lane1;
  assign execute_ctrl2_down_Decode_UOP_ID_lane1 = execute_ctrl2_up_Decode_UOP_ID_lane1;
  assign execute_ctrl2_down_RS1_RFID_lane1 = execute_ctrl2_up_RS1_RFID_lane1;
  assign execute_ctrl2_down_RS1_PHYS_lane1 = execute_ctrl2_up_RS1_PHYS_lane1;
  assign execute_ctrl2_down_RS2_RFID_lane1 = execute_ctrl2_up_RS2_RFID_lane1;
  assign execute_ctrl2_down_RS2_PHYS_lane1 = execute_ctrl2_up_RS2_PHYS_lane1;
  assign execute_ctrl2_down_RD_RFID_lane1 = execute_ctrl2_up_RD_RFID_lane1;
  assign execute_ctrl2_down_RD_PHYS_lane1 = execute_ctrl2_up_RD_PHYS_lane1;
  assign execute_ctrl2_down_LANE_AGE_lane1 = execute_ctrl2_up_LANE_AGE_lane1;
  assign execute_ctrl2_down_AguPlugin_SIZE_lane0 = execute_ctrl2_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  assign execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 = execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1;
  assign execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1 = execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1;
  assign execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0 = execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  assign execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1 = execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1;
  assign execute_ctrl2_down_float_RS1_lane0 = execute_ctrl2_up_float_RS1_lane0;
  assign execute_ctrl2_down_float_RS2_lane0 = execute_ctrl2_up_float_RS2_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_SEL_lane0 = execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_DivPlugin_SEL_lane0 = execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_SEL_lane0 = execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  assign execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0 = execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl2_down_late0_BranchPlugin_SEL_lane0 = execute_ctrl2_up_late0_BranchPlugin_SEL_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuCsrPlugin_DIRTY_lane0 = execute_ctrl2_up_FpuCsrPlugin_DIRTY_lane0;
  assign execute_ctrl2_down_FpuClassPlugin_SEL_lane0 = execute_ctrl2_up_FpuClassPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_SEL_FLOAT_lane0 = execute_ctrl2_up_FpuCmpPlugin_SEL_FLOAT_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_SEL_CMP_lane0 = execute_ctrl2_up_FpuCmpPlugin_SEL_CMP_lane0;
  assign execute_ctrl2_down_FpuF2iPlugin_SEL_lane0 = execute_ctrl2_up_FpuF2iPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuMvPlugin_SEL_FLOAT_lane0 = execute_ctrl2_up_FpuMvPlugin_SEL_FLOAT_lane0;
  assign execute_ctrl2_down_FpuMvPlugin_SEL_INT_lane0 = execute_ctrl2_up_FpuMvPlugin_SEL_INT_lane0;
  assign execute_ctrl2_down_AguPlugin_SEL_lane0 = execute_ctrl2_up_AguPlugin_SEL_lane0;
  assign execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl2_down_FpuAddPlugin_SEL_lane0 = execute_ctrl2_up_FpuAddPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuMulPlugin_SEL_lane0 = execute_ctrl2_up_FpuMulPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuSqrtPlugin_SEL_lane0 = execute_ctrl2_up_FpuSqrtPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuXxPlugin_SEL_lane0 = execute_ctrl2_up_FpuXxPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuDivPlugin_SEL_lane0 = execute_ctrl2_up_FpuDivPlugin_SEL_lane0;
  assign execute_ctrl2_down_FpuUnpackerPlugin_SEL_I2F_lane0 = execute_ctrl2_up_FpuUnpackerPlugin_SEL_I2F_lane0;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl2_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl2_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_4_lane0 = execute_ctrl2_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_7_lane0 = execute_ctrl2_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_11_lane0 = execute_ctrl2_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_3_lane0 = execute_ctrl2_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_5_lane0 = execute_ctrl2_up_COMPLETION_AT_5_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_8_lane0 = execute_ctrl2_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_2_lane0 = execute_ctrl2_up_COMPLETION_AT_2_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl2_down_SrcStageables_REVERT_lane0 = execute_ctrl2_up_SrcStageables_REVERT_lane0;
  assign execute_ctrl2_down_SrcStageables_ZERO_lane0 = execute_ctrl2_up_SrcStageables_ZERO_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_3_lane0 = execute_ctrl2_up_BYPASSED_AT_3_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_4_lane0 = execute_ctrl2_up_BYPASSED_AT_4_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_5_lane0 = execute_ctrl2_up_BYPASSED_AT_5_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_6_lane0 = execute_ctrl2_up_BYPASSED_AT_6_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_7_lane0 = execute_ctrl2_up_BYPASSED_AT_7_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_8_lane0 = execute_ctrl2_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_9_lane0 = execute_ctrl2_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_10_lane0 = execute_ctrl2_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 = execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 = execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 = execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  assign execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl2_down_MulPlugin_HIGH_lane0 = execute_ctrl2_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  assign execute_ctrl2_down_DivPlugin_REM_lane0 = execute_ctrl2_up_DivPlugin_REM_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign execute_ctrl2_down_FpuUtils_FORMAT_lane0 = execute_ctrl2_up_FpuUtils_FORMAT_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0 = execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_INVERT_lane0 = execute_ctrl2_up_FpuCmpPlugin_INVERT_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_SGNJ_RS1_lane0 = execute_ctrl2_up_FpuCmpPlugin_SGNJ_RS1_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_LESS_lane0 = execute_ctrl2_up_FpuCmpPlugin_LESS_lane0;
  assign execute_ctrl2_down_FpuCmpPlugin_EQUAL_lane0 = execute_ctrl2_up_FpuCmpPlugin_EQUAL_lane0;
  assign execute_ctrl2_down_AguPlugin_LOAD_lane0 = execute_ctrl2_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl2_down_AguPlugin_STORE_lane0 = execute_ctrl2_up_AguPlugin_STORE_lane0;
  assign execute_ctrl2_down_AguPlugin_ATOMIC_lane0 = execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl2_down_AguPlugin_FLOAT_lane0 = execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_OP_lane0 = execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  assign execute_ctrl2_down_FpuAddPlugin_SUB_lane0 = execute_ctrl2_up_FpuAddPlugin_SUB_lane0;
  assign execute_ctrl2_down_FpuMulPlugin_FMA_lane0 = execute_ctrl2_up_FpuMulPlugin_FMA_lane0;
  assign execute_ctrl2_down_FpuMulPlugin_SUB1_lane0 = execute_ctrl2_up_FpuMulPlugin_SUB1_lane0;
  assign execute_ctrl2_down_FpuMulPlugin_SUB2_lane0 = execute_ctrl2_up_FpuMulPlugin_SUB2_lane0;
  assign execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  assign execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  assign execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1 = execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1;
  assign execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1 = execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1;
  assign execute_ctrl2_down_early1_BranchPlugin_SEL_lane1 = execute_ctrl2_up_early1_BranchPlugin_SEL_lane1;
  assign execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1 = execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1;
  assign execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1 = execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign execute_ctrl2_down_late1_BranchPlugin_SEL_lane1 = execute_ctrl2_up_late1_BranchPlugin_SEL_lane1;
  assign execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1 = execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign execute_ctrl2_down_COMPLETION_AT_2_lane1 = execute_ctrl2_up_COMPLETION_AT_2_lane1;
  assign execute_ctrl2_down_COMPLETION_AT_4_lane1 = execute_ctrl2_up_COMPLETION_AT_4_lane1;
  assign execute_ctrl2_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = execute_ctrl2_up_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  assign execute_ctrl2_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = execute_ctrl2_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  assign execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1 = execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1;
  assign execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign execute_ctrl2_down_SrcStageables_REVERT_lane1 = execute_ctrl2_up_SrcStageables_REVERT_lane1;
  assign execute_ctrl2_down_SrcStageables_ZERO_lane1 = execute_ctrl2_up_SrcStageables_ZERO_lane1;
  assign execute_ctrl2_down_BYPASSED_AT_3_lane1 = execute_ctrl2_up_BYPASSED_AT_3_lane1;
  assign execute_ctrl2_down_SrcStageables_UNSIGNED_lane1 = execute_ctrl2_up_SrcStageables_UNSIGNED_lane1;
  assign execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 = execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1;
  assign execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1 = execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1;
  assign execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 = execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1 = execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  assign execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  assign execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX = execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  assign execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF = execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  assign execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF = execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  assign execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ = execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  assign execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV = execute_ctrl2_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  assign execute_ctrl2_down_COMMIT_lane1 = execute_ctrl2_up_COMMIT_lane1;
  assign execute_ctrl3_up_ready = execute_ctrl3_down_isReady;
  assign execute_ctrl3_down_Decode_UOP_lane0 = execute_ctrl3_up_Decode_UOP_lane0;
  assign execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  assign execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl3_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 = execute_ctrl3_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
  assign execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl3_down_PC_lane0 = execute_ctrl3_up_PC_lane0;
  assign execute_ctrl3_down_TRAP_lane0 = execute_ctrl3_up_TRAP_lane0;
  assign execute_ctrl3_down_Decode_UOP_ID_lane0 = execute_ctrl3_up_Decode_UOP_ID_lane0;
  assign execute_ctrl3_down_RS1_RFID_lane0 = execute_ctrl3_up_RS1_RFID_lane0;
  assign execute_ctrl3_down_RS1_PHYS_lane0 = execute_ctrl3_up_RS1_PHYS_lane0;
  assign execute_ctrl3_down_RS2_RFID_lane0 = execute_ctrl3_up_RS2_RFID_lane0;
  assign execute_ctrl3_down_RS2_PHYS_lane0 = execute_ctrl3_up_RS2_PHYS_lane0;
  assign execute_ctrl3_down_RD_RFID_lane0 = execute_ctrl3_up_RD_RFID_lane0;
  assign execute_ctrl3_down_RD_PHYS_lane0 = execute_ctrl3_up_RD_PHYS_lane0;
  assign execute_ctrl3_down_LANE_AGE_lane0 = execute_ctrl3_up_LANE_AGE_lane0;
  assign execute_ctrl3_down_Decode_UOP_lane1 = execute_ctrl3_up_Decode_UOP_lane1;
  assign execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1 = execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1;
  assign execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1 = execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1 = execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1;
  assign execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign execute_ctrl3_down_PC_lane1 = execute_ctrl3_up_PC_lane1;
  assign execute_ctrl3_down_TRAP_lane1 = execute_ctrl3_up_TRAP_lane1;
  assign execute_ctrl3_down_Decode_UOP_ID_lane1 = execute_ctrl3_up_Decode_UOP_ID_lane1;
  assign execute_ctrl3_down_RS1_RFID_lane1 = execute_ctrl3_up_RS1_RFID_lane1;
  assign execute_ctrl3_down_RS1_PHYS_lane1 = execute_ctrl3_up_RS1_PHYS_lane1;
  assign execute_ctrl3_down_RS2_RFID_lane1 = execute_ctrl3_up_RS2_RFID_lane1;
  assign execute_ctrl3_down_RS2_PHYS_lane1 = execute_ctrl3_up_RS2_PHYS_lane1;
  assign execute_ctrl3_down_RD_RFID_lane1 = execute_ctrl3_up_RD_RFID_lane1;
  assign execute_ctrl3_down_RD_PHYS_lane1 = execute_ctrl3_up_RD_PHYS_lane1;
  assign execute_ctrl3_down_LANE_AGE_lane1 = execute_ctrl3_up_LANE_AGE_lane1;
  assign execute_ctrl3_down_COMPLETED_lane1 = execute_ctrl3_up_COMPLETED_lane1;
  assign execute_ctrl3_down_AguPlugin_SIZE_lane0 = execute_ctrl3_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl3_down_float_RS2_lane0 = execute_ctrl3_up_float_RS2_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_SEL_lane0 = execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl3_down_early0_DivPlugin_SEL_lane0 = execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0 = execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl3_down_late0_BranchPlugin_SEL_lane0 = execute_ctrl3_up_late0_BranchPlugin_SEL_lane0;
  assign execute_ctrl3_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl3_down_FpuCsrPlugin_DIRTY_lane0 = execute_ctrl3_up_FpuCsrPlugin_DIRTY_lane0;
  assign execute_ctrl3_down_FpuClassPlugin_SEL_lane0 = execute_ctrl3_up_FpuClassPlugin_SEL_lane0;
  assign execute_ctrl3_down_FpuCmpPlugin_SEL_FLOAT_lane0 = execute_ctrl3_up_FpuCmpPlugin_SEL_FLOAT_lane0;
  assign execute_ctrl3_down_FpuCmpPlugin_SEL_CMP_lane0 = execute_ctrl3_up_FpuCmpPlugin_SEL_CMP_lane0;
  assign execute_ctrl3_down_FpuF2iPlugin_SEL_lane0 = execute_ctrl3_up_FpuF2iPlugin_SEL_lane0;
  assign execute_ctrl3_down_FpuMvPlugin_SEL_FLOAT_lane0 = execute_ctrl3_up_FpuMvPlugin_SEL_FLOAT_lane0;
  assign execute_ctrl3_down_FpuMvPlugin_SEL_INT_lane0 = execute_ctrl3_up_FpuMvPlugin_SEL_INT_lane0;
  assign execute_ctrl3_down_AguPlugin_SEL_lane0 = execute_ctrl3_up_AguPlugin_SEL_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_SEL_lane0 = execute_ctrl3_up_FpuMulPlugin_SEL_lane0;
  assign execute_ctrl3_down_FpuXxPlugin_SEL_lane0 = execute_ctrl3_up_FpuXxPlugin_SEL_lane0;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl3_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl3_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_4_lane0 = execute_ctrl3_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_7_lane0 = execute_ctrl3_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_11_lane0 = execute_ctrl3_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_3_lane0 = execute_ctrl3_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_5_lane0 = execute_ctrl3_up_COMPLETION_AT_5_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_8_lane0 = execute_ctrl3_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl3_down_SrcStageables_REVERT_lane0 = execute_ctrl3_up_SrcStageables_REVERT_lane0;
  assign execute_ctrl3_down_SrcStageables_ZERO_lane0 = execute_ctrl3_up_SrcStageables_ZERO_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_4_lane0 = execute_ctrl3_up_BYPASSED_AT_4_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_5_lane0 = execute_ctrl3_up_BYPASSED_AT_5_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_6_lane0 = execute_ctrl3_up_BYPASSED_AT_6_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_7_lane0 = execute_ctrl3_up_BYPASSED_AT_7_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_8_lane0 = execute_ctrl3_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_9_lane0 = execute_ctrl3_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl3_down_BYPASSED_AT_10_lane0 = execute_ctrl3_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl3_down_SrcStageables_UNSIGNED_lane0 = execute_ctrl3_up_SrcStageables_UNSIGNED_lane0;
  assign execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0 = execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0;
  assign execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0 = execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0;
  assign execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl3_down_MulPlugin_HIGH_lane0 = execute_ctrl3_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl3_down_FpuUtils_FORMAT_lane0 = execute_ctrl3_up_FpuUtils_FORMAT_lane0;
  assign execute_ctrl3_down_FpuCmpPlugin_FLOAT_OP_lane0 = execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0;
  assign execute_ctrl3_down_AguPlugin_LOAD_lane0 = execute_ctrl3_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl3_down_AguPlugin_STORE_lane0 = execute_ctrl3_up_AguPlugin_STORE_lane0;
  assign execute_ctrl3_down_AguPlugin_ATOMIC_lane0 = execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl3_down_AguPlugin_FLOAT_lane0 = execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_FMA_lane0 = execute_ctrl3_up_FpuMulPlugin_FMA_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_SUB1_lane0 = execute_ctrl3_up_FpuMulPlugin_SUB1_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_SUB2_lane0 = execute_ctrl3_up_FpuMulPlugin_SUB2_lane0;
  assign execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  assign execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  assign execute_ctrl3_down_early1_BranchPlugin_SEL_lane1 = execute_ctrl3_up_early1_BranchPlugin_SEL_lane1;
  assign execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1 = execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1;
  assign execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1 = execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign execute_ctrl3_down_late1_BranchPlugin_SEL_lane1 = execute_ctrl3_up_late1_BranchPlugin_SEL_lane1;
  assign execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1 = execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign execute_ctrl3_down_COMPLETION_AT_4_lane1 = execute_ctrl3_up_COMPLETION_AT_4_lane1;
  assign execute_ctrl3_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = execute_ctrl3_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  assign execute_ctrl3_down_SrcStageables_REVERT_lane1 = execute_ctrl3_up_SrcStageables_REVERT_lane1;
  assign execute_ctrl3_down_SrcStageables_ZERO_lane1 = execute_ctrl3_up_SrcStageables_ZERO_lane1;
  assign execute_ctrl3_down_SrcStageables_UNSIGNED_lane1 = execute_ctrl3_up_SrcStageables_UNSIGNED_lane1;
  assign execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1 = execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1;
  assign execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1 = execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1;
  assign execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1 = execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1 = execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  assign execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  assign execute_ctrl3_down_COMMIT_lane0 = execute_ctrl3_up_COMMIT_lane0;
  assign execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX = execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
  assign execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF = execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
  assign execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF = execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
  assign execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ = execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
  assign execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV = execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
  assign execute_ctrl3_down_COMMIT_lane1 = execute_ctrl3_up_COMMIT_lane1;
  assign execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0 = execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  assign execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  assign execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0 = execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign execute_ctrl3_down_FpuUtils_ROUNDING_lane0 = execute_ctrl3_up_FpuUtils_ROUNDING_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_WB_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_WB_lane0;
  assign execute_ctrl3_down_LsuL1_MASK_lane0 = execute_ctrl3_up_LsuL1_MASK_lane0;
  assign execute_ctrl3_down_LsuL1_SIZE_lane0 = execute_ctrl3_up_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuL1_LOAD_lane0 = execute_ctrl3_up_LsuL1_LOAD_lane0;
  assign execute_ctrl3_down_LsuL1_ATOMIC_lane0 = execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl3_down_LsuL1_STORE_lane0 = execute_ctrl3_up_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuL1_CLEAN_lane0 = execute_ctrl3_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl3_down_LsuL1_INVALID_lane0 = execute_ctrl3_up_LsuL1_INVALID_lane0;
  assign execute_ctrl3_down_LsuL1_PREFETCH_lane0 = execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl3_down_LsuL1_FLUSH_lane0 = execute_ctrl3_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl3_down_Decode_STORE_ID_lane0 = execute_ctrl3_up_Decode_STORE_ID_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl3_down_LsuPlugin_SB_PTR_lane0 = execute_ctrl3_up_LsuPlugin_SB_PTR_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0 = execute_ctrl3_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0 = execute_ctrl3_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  assign execute_ctrl3_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0 = execute_ctrl3_up_FpuUnpack_RS1_IS_SUBNORMAL_lane0;
  assign execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode = execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode;
  assign execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet = execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_quiet;
  assign execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign = execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_sign;
  assign execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent = _zz_execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mantissa = execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mantissa;
  assign execute_ctrl3_down_FpuUnpack_RS1_badBoxing_HIT_lane0 = execute_ctrl3_up_FpuUnpack_RS1_badBoxing_HIT_lane0;
  assign execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode = execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode;
  assign execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_quiet = execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_quiet;
  assign execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_sign = execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_sign;
  assign execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent = _zz_execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mantissa = execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mantissa;
  assign execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode = execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode;
  assign execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_quiet = execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_quiet;
  assign execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_sign = execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_sign;
  assign execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent = _zz_execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mantissa = execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mantissa;
  assign execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  assign execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0 = execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0;
  assign execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0 = execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
  assign execute_ctrl3_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0 = execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
  assign execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 = execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
  assign execute_ctrl3_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 = execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = _zz_execute_ctrl3_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_SIGN_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  assign execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 = execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  assign execute_ctrl4_up_ready = execute_ctrl4_down_isReady;
  assign execute_ctrl4_down_Decode_UOP_lane0 = execute_ctrl4_up_Decode_UOP_lane0;
  assign execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 = execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
  assign execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl4_down_PC_lane0 = execute_ctrl4_up_PC_lane0;
  assign execute_ctrl4_down_Decode_UOP_ID_lane0 = execute_ctrl4_up_Decode_UOP_ID_lane0;
  assign execute_ctrl4_down_RD_RFID_lane0 = execute_ctrl4_up_RD_RFID_lane0;
  assign execute_ctrl4_down_RD_PHYS_lane0 = execute_ctrl4_up_RD_PHYS_lane0;
  assign execute_ctrl4_down_LANE_AGE_lane0 = execute_ctrl4_up_LANE_AGE_lane0;
  assign execute_ctrl4_down_Decode_UOP_lane1 = execute_ctrl4_up_Decode_UOP_lane1;
  assign execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1 = execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1;
  assign execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1 = execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1 = execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1;
  assign execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign execute_ctrl4_down_PC_lane1 = execute_ctrl4_up_PC_lane1;
  assign execute_ctrl4_down_TRAP_lane1 = execute_ctrl4_up_TRAP_lane1;
  assign execute_ctrl4_down_Decode_UOP_ID_lane1 = execute_ctrl4_up_Decode_UOP_ID_lane1;
  assign execute_ctrl4_down_RD_RFID_lane1 = execute_ctrl4_up_RD_RFID_lane1;
  assign execute_ctrl4_down_RD_PHYS_lane1 = execute_ctrl4_up_RD_PHYS_lane1;
  assign execute_ctrl4_down_LANE_AGE_lane1 = execute_ctrl4_up_LANE_AGE_lane1;
  assign execute_ctrl4_down_AguPlugin_SIZE_lane0 = execute_ctrl4_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl4_down_integer_RS2_lane0 = execute_ctrl4_up_integer_RS2_lane0;
  assign execute_ctrl4_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl4_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_SEL_lane0 = execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0 = execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl4_down_late0_BranchPlugin_SEL_lane0 = execute_ctrl4_up_late0_BranchPlugin_SEL_lane0;
  assign execute_ctrl4_down_FpuCsrPlugin_DIRTY_lane0 = execute_ctrl4_up_FpuCsrPlugin_DIRTY_lane0;
  assign execute_ctrl4_down_FpuF2iPlugin_SEL_lane0 = execute_ctrl4_up_FpuF2iPlugin_SEL_lane0;
  assign execute_ctrl4_down_FpuMvPlugin_SEL_FLOAT_lane0 = execute_ctrl4_up_FpuMvPlugin_SEL_FLOAT_lane0;
  assign execute_ctrl4_down_AguPlugin_SEL_lane0 = execute_ctrl4_up_AguPlugin_SEL_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_SEL_lane0 = execute_ctrl4_up_FpuMulPlugin_SEL_lane0;
  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl4_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl4_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_4_lane0 = execute_ctrl4_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_7_lane0 = execute_ctrl4_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_11_lane0 = execute_ctrl4_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_5_lane0 = execute_ctrl4_up_COMPLETION_AT_5_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_8_lane0 = execute_ctrl4_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl4_down_SrcStageables_REVERT_lane0 = execute_ctrl4_up_SrcStageables_REVERT_lane0;
  assign execute_ctrl4_down_SrcStageables_ZERO_lane0 = execute_ctrl4_up_SrcStageables_ZERO_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_5_lane0 = execute_ctrl4_up_BYPASSED_AT_5_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_6_lane0 = execute_ctrl4_up_BYPASSED_AT_6_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_7_lane0 = execute_ctrl4_up_BYPASSED_AT_7_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_8_lane0 = execute_ctrl4_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_9_lane0 = execute_ctrl4_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl4_down_BYPASSED_AT_10_lane0 = execute_ctrl4_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl4_down_SrcStageables_UNSIGNED_lane0 = execute_ctrl4_up_SrcStageables_UNSIGNED_lane0;
  assign execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 = execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0;
  assign execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0 = execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0;
  assign execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl4_down_MulPlugin_HIGH_lane0 = execute_ctrl4_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl4_down_FpuUtils_FORMAT_lane0 = execute_ctrl4_up_FpuUtils_FORMAT_lane0;
  assign execute_ctrl4_down_AguPlugin_LOAD_lane0 = execute_ctrl4_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl4_down_AguPlugin_STORE_lane0 = execute_ctrl4_up_AguPlugin_STORE_lane0;
  assign execute_ctrl4_down_AguPlugin_ATOMIC_lane0 = execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl4_down_AguPlugin_FLOAT_lane0 = execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_FMA_lane0 = execute_ctrl4_up_FpuMulPlugin_FMA_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_SUB1_lane0 = execute_ctrl4_up_FpuMulPlugin_SUB1_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_SUB2_lane0 = execute_ctrl4_up_FpuMulPlugin_SUB2_lane0;
  assign execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl4_down_early1_BranchPlugin_SEL_lane1 = execute_ctrl4_up_early1_BranchPlugin_SEL_lane1;
  assign execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1 = execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1;
  assign execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1 = execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign execute_ctrl4_down_late1_BranchPlugin_SEL_lane1 = execute_ctrl4_up_late1_BranchPlugin_SEL_lane1;
  assign execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1 = execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign execute_ctrl4_down_COMPLETION_AT_4_lane1 = execute_ctrl4_up_COMPLETION_AT_4_lane1;
  assign execute_ctrl4_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = execute_ctrl4_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  assign execute_ctrl4_down_SrcStageables_REVERT_lane1 = execute_ctrl4_up_SrcStageables_REVERT_lane1;
  assign execute_ctrl4_down_SrcStageables_ZERO_lane1 = execute_ctrl4_up_SrcStageables_ZERO_lane1;
  assign execute_ctrl4_down_SrcStageables_UNSIGNED_lane1 = execute_ctrl4_up_SrcStageables_UNSIGNED_lane1;
  assign execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 = execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1;
  assign execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1 = execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1;
  assign execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 = execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1 = execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign execute_ctrl4_down_COMMIT_lane1 = execute_ctrl4_up_COMMIT_lane1;
  assign execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_4_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_5_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_6_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_7_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_8_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_9_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_10_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_11_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_12_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_13_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_14_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_15_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0;
  assign execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign execute_ctrl4_down_FpuUtils_ROUNDING_lane0 = execute_ctrl4_up_FpuUtils_ROUNDING_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_WB_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_WB_lane0;
  assign execute_ctrl4_down_LsuL1_MASK_lane0 = execute_ctrl4_up_LsuL1_MASK_lane0;
  assign execute_ctrl4_down_LsuL1_SIZE_lane0 = execute_ctrl4_up_LsuL1_SIZE_lane0;
  assign execute_ctrl4_down_LsuL1_LOAD_lane0 = execute_ctrl4_up_LsuL1_LOAD_lane0;
  assign execute_ctrl4_down_LsuL1_ATOMIC_lane0 = execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl4_down_LsuL1_STORE_lane0 = execute_ctrl4_up_LsuL1_STORE_lane0;
  assign execute_ctrl4_down_LsuL1_CLEAN_lane0 = execute_ctrl4_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl4_down_LsuL1_INVALID_lane0 = execute_ctrl4_up_LsuL1_INVALID_lane0;
  assign execute_ctrl4_down_LsuL1_PREFETCH_lane0 = execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuL1_FLUSH_lane0 = execute_ctrl4_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl4_down_Decode_STORE_ID_lane0 = execute_ctrl4_up_Decode_STORE_ID_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuPlugin_SB_PTR_lane0 = execute_ctrl4_up_LsuPlugin_SB_PTR_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0 = execute_ctrl4_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0 = execute_ctrl4_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
  assign execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode = execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode;
  assign execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_quiet = execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_quiet;
  assign execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign = execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_sign;
  assign execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent = _zz_execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mantissa = execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mantissa;
  assign execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode = execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode;
  assign execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_quiet = execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_quiet;
  assign execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_sign = execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_sign;
  assign execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent = _zz_execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mantissa = execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mantissa;
  assign execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode = execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode;
  assign execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_quiet = execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_quiet;
  assign execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_sign = execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_sign;
  assign execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent = _zz_execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mantissa = execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mantissa;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = _zz_execute_ctrl4_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_SIGN_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  assign execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 = execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  assign execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  assign execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 = execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0;
  assign execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0 = execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0;
  assign execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 = execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1;
  assign execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1 = execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_2_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  assign execute_ctrl4_down_MMU_TRANSLATED_lane0 = execute_ctrl4_up_MMU_TRANSLATED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  assign execute_ctrl4_down_MMU_ACCESS_FAULT_lane0 = execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  assign execute_ctrl4_down_MMU_REFILL_lane0 = execute_ctrl4_up_MMU_REFILL_lane0;
  assign execute_ctrl4_down_MMU_HAZARD_lane0 = execute_ctrl4_up_MMU_HAZARD_lane0;
  assign execute_ctrl4_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 = execute_ctrl4_up_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
  assign execute_ctrl4_down_FpuF2iPlugin_logic_onShift_resign_lane0 = execute_ctrl4_up_FpuF2iPlugin_logic_onShift_resign_lane0;
  assign execute_ctrl4_down_FpuF2iPlugin_logic_onShift_increment_lane0 = execute_ctrl4_up_FpuF2iPlugin_logic_onShift_increment_lane0;
  assign execute_ctrl4_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0 = execute_ctrl4_up_FpuF2iPlugin_logic_onShift_incrementPatched_lane0;
  assign execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0 = execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  assign execute_ctrl5_up_ready = execute_ctrl5_down_isReady;
  assign execute_ctrl5_down_LANE_SEL_lane0 = execute_ctrl5_up_LANE_SEL_lane0;
  assign execute_ctrl5_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl5_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl5_down_TRAP_lane0 = execute_ctrl5_up_TRAP_lane0;
  assign execute_ctrl5_down_Decode_UOP_ID_lane0 = execute_ctrl5_up_Decode_UOP_ID_lane0;
  assign execute_ctrl5_down_RD_ENABLE_lane0 = execute_ctrl5_up_RD_ENABLE_lane0;
  assign execute_ctrl5_down_RD_RFID_lane0 = execute_ctrl5_up_RD_RFID_lane0;
  assign execute_ctrl5_down_RD_PHYS_lane0 = execute_ctrl5_up_RD_PHYS_lane0;
  assign execute_ctrl5_down_LANE_AGE_lane0 = execute_ctrl5_up_LANE_AGE_lane0;
  assign execute_ctrl5_down_LANE_SEL_lane1 = execute_ctrl5_up_LANE_SEL_lane1;
  assign execute_ctrl5_down_RD_RFID_lane1 = execute_ctrl5_up_RD_RFID_lane1;
  assign execute_ctrl5_down_RD_PHYS_lane1 = execute_ctrl5_up_RD_PHYS_lane1;
  assign execute_ctrl5_down_LANE_AGE_lane1 = execute_ctrl5_up_LANE_AGE_lane1;
  assign execute_ctrl5_down_FpuMulPlugin_SEL_lane0 = execute_ctrl5_up_FpuMulPlugin_SEL_lane0;
  assign execute_ctrl5_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl5_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl5_down_COMPLETION_AT_7_lane0 = execute_ctrl5_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl5_down_COMPLETION_AT_11_lane0 = execute_ctrl5_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl5_down_COMPLETION_AT_5_lane0 = execute_ctrl5_up_COMPLETION_AT_5_lane0;
  assign execute_ctrl5_down_COMPLETION_AT_8_lane0 = execute_ctrl5_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl5_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl5_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl5_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl5_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl5_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0 = execute_ctrl5_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
  assign execute_ctrl5_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl5_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl5_down_BYPASSED_AT_6_lane0 = execute_ctrl5_up_BYPASSED_AT_6_lane0;
  assign execute_ctrl5_down_BYPASSED_AT_7_lane0 = execute_ctrl5_up_BYPASSED_AT_7_lane0;
  assign execute_ctrl5_down_BYPASSED_AT_8_lane0 = execute_ctrl5_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl5_down_BYPASSED_AT_9_lane0 = execute_ctrl5_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl5_down_BYPASSED_AT_10_lane0 = execute_ctrl5_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl5_down_FpuUtils_FORMAT_lane0 = execute_ctrl5_up_FpuUtils_FORMAT_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_FMA_lane0 = execute_ctrl5_up_FpuMulPlugin_FMA_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_SUB1_lane0 = execute_ctrl5_up_FpuMulPlugin_SUB1_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_SUB2_lane0 = execute_ctrl5_up_FpuMulPlugin_SUB2_lane0;
  assign execute_ctrl5_down_COMMIT_lane0 = execute_ctrl5_up_COMMIT_lane0;
  assign execute_ctrl5_down_COMMIT_lane1 = execute_ctrl5_up_COMMIT_lane1;
  assign execute_ctrl5_down_FpuUtils_ROUNDING_lane0 = execute_ctrl5_up_FpuUtils_ROUNDING_lane0;
  assign execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mode = execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode;
  assign execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_quiet = execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_quiet;
  assign execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_sign = execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_sign;
  assign execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_exponent = _zz_execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_exponent;
  assign execute_ctrl5_down_FpuUnpack_RS1_RS_lane0_mantissa = execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mantissa;
  assign execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mode = execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode;
  assign execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_quiet = execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_quiet;
  assign execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_sign = execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_sign;
  assign execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_exponent = _zz_execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_exponent;
  assign execute_ctrl5_down_FpuUnpack_RS2_RS_lane0_mantissa = execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mantissa;
  assign execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mode = execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode;
  assign execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_quiet = execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_quiet;
  assign execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_sign = execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_sign;
  assign execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent = _zz_execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_exponent;
  assign execute_ctrl5_down_FpuUnpack_RS3_RS_lane0_mantissa = execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mantissa;
  assign execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0 = _zz_execute_ctrl5_down_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_SIGN_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_SIGN_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
  assign execute_ctrl5_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0 = execute_ctrl5_up_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
  assign execute_ctrl6_up_ready = execute_ctrl6_down_isReady;
  assign execute_ctrl6_down_LANE_SEL_lane0 = execute_ctrl6_up_LANE_SEL_lane0;
  assign execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl6_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl6_down_TRAP_lane0 = execute_ctrl6_up_TRAP_lane0;
  assign execute_ctrl6_down_Decode_UOP_ID_lane0 = execute_ctrl6_up_Decode_UOP_ID_lane0;
  assign execute_ctrl6_down_RD_ENABLE_lane0 = execute_ctrl6_up_RD_ENABLE_lane0;
  assign execute_ctrl6_down_RD_RFID_lane0 = execute_ctrl6_up_RD_RFID_lane0;
  assign execute_ctrl6_down_RD_PHYS_lane0 = execute_ctrl6_up_RD_PHYS_lane0;
  assign execute_ctrl6_down_LANE_AGE_lane0 = execute_ctrl6_up_LANE_AGE_lane0;
  assign execute_ctrl6_down_COMPLETED_lane0 = execute_ctrl6_up_COMPLETED_lane0;
  assign execute_ctrl6_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl6_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl6_down_COMPLETION_AT_7_lane0 = execute_ctrl6_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl6_down_COMPLETION_AT_11_lane0 = execute_ctrl6_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl6_down_COMPLETION_AT_8_lane0 = execute_ctrl6_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl6_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl6_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl6_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl6_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl6_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl6_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl6_down_BYPASSED_AT_7_lane0 = execute_ctrl6_up_BYPASSED_AT_7_lane0;
  assign execute_ctrl6_down_BYPASSED_AT_8_lane0 = execute_ctrl6_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl6_down_BYPASSED_AT_9_lane0 = execute_ctrl6_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl6_down_BYPASSED_AT_10_lane0 = execute_ctrl6_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl6_down_COMMIT_lane0 = execute_ctrl6_up_COMMIT_lane0;
  assign execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl6_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  assign execute_ctrl7_up_ready = execute_ctrl7_down_isReady;
  assign execute_ctrl7_down_LANE_SEL_lane0 = execute_ctrl7_up_LANE_SEL_lane0;
  assign execute_ctrl7_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 = execute_ctrl7_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
  assign execute_ctrl7_down_TRAP_lane0 = execute_ctrl7_up_TRAP_lane0;
  assign execute_ctrl7_down_Decode_UOP_ID_lane0 = execute_ctrl7_up_Decode_UOP_ID_lane0;
  assign execute_ctrl7_down_RD_ENABLE_lane0 = execute_ctrl7_up_RD_ENABLE_lane0;
  assign execute_ctrl7_down_RD_RFID_lane0 = execute_ctrl7_up_RD_RFID_lane0;
  assign execute_ctrl7_down_RD_PHYS_lane0 = execute_ctrl7_up_RD_PHYS_lane0;
  assign execute_ctrl7_down_LANE_AGE_lane0 = execute_ctrl7_up_LANE_AGE_lane0;
  assign execute_ctrl7_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl7_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl7_down_COMPLETION_AT_7_lane0 = execute_ctrl7_up_COMPLETION_AT_7_lane0;
  assign execute_ctrl7_down_COMPLETION_AT_11_lane0 = execute_ctrl7_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl7_down_COMPLETION_AT_8_lane0 = execute_ctrl7_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl7_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl7_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl7_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl7_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl7_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl7_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl7_down_BYPASSED_AT_8_lane0 = execute_ctrl7_up_BYPASSED_AT_8_lane0;
  assign execute_ctrl7_down_BYPASSED_AT_9_lane0 = execute_ctrl7_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl7_down_BYPASSED_AT_10_lane0 = execute_ctrl7_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl7_down_COMMIT_lane0 = execute_ctrl7_up_COMMIT_lane0;
  assign execute_ctrl8_up_ready = execute_ctrl8_down_isReady;
  assign execute_ctrl8_down_LANE_SEL_lane0 = execute_ctrl8_up_LANE_SEL_lane0;
  assign execute_ctrl8_down_TRAP_lane0 = execute_ctrl8_up_TRAP_lane0;
  assign execute_ctrl8_down_Decode_UOP_ID_lane0 = execute_ctrl8_up_Decode_UOP_ID_lane0;
  assign execute_ctrl8_down_RD_ENABLE_lane0 = execute_ctrl8_up_RD_ENABLE_lane0;
  assign execute_ctrl8_down_RD_RFID_lane0 = execute_ctrl8_up_RD_RFID_lane0;
  assign execute_ctrl8_down_RD_PHYS_lane0 = execute_ctrl8_up_RD_PHYS_lane0;
  assign execute_ctrl8_down_LANE_AGE_lane0 = execute_ctrl8_up_LANE_AGE_lane0;
  assign execute_ctrl8_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl8_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl8_down_COMPLETION_AT_11_lane0 = execute_ctrl8_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl8_down_COMPLETION_AT_8_lane0 = execute_ctrl8_up_COMPLETION_AT_8_lane0;
  assign execute_ctrl8_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl8_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl8_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0 = execute_ctrl8_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
  assign execute_ctrl8_down_BYPASSED_AT_9_lane0 = execute_ctrl8_up_BYPASSED_AT_9_lane0;
  assign execute_ctrl8_down_BYPASSED_AT_10_lane0 = execute_ctrl8_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl8_down_COMMIT_lane0 = execute_ctrl8_up_COMMIT_lane0;
  assign execute_ctrl9_up_ready = execute_ctrl9_down_isReady;
  assign execute_ctrl9_down_LANE_SEL_lane0 = execute_ctrl9_up_LANE_SEL_lane0;
  assign execute_ctrl9_down_TRAP_lane0 = execute_ctrl9_up_TRAP_lane0;
  assign execute_ctrl9_down_Decode_UOP_ID_lane0 = execute_ctrl9_up_Decode_UOP_ID_lane0;
  assign execute_ctrl9_down_RD_ENABLE_lane0 = execute_ctrl9_up_RD_ENABLE_lane0;
  assign execute_ctrl9_down_RD_RFID_lane0 = execute_ctrl9_up_RD_RFID_lane0;
  assign execute_ctrl9_down_RD_PHYS_lane0 = execute_ctrl9_up_RD_PHYS_lane0;
  assign execute_ctrl9_down_LANE_AGE_lane0 = execute_ctrl9_up_LANE_AGE_lane0;
  assign execute_ctrl9_down_COMPLETED_lane0 = execute_ctrl9_up_COMPLETED_lane0;
  assign execute_ctrl9_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl9_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl9_down_COMPLETION_AT_11_lane0 = execute_ctrl9_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl9_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl9_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl9_down_BYPASSED_AT_10_lane0 = execute_ctrl9_up_BYPASSED_AT_10_lane0;
  assign execute_ctrl9_down_COMMIT_lane0 = execute_ctrl9_up_COMMIT_lane0;
  assign execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl9_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  assign execute_ctrl10_up_ready = execute_ctrl10_down_isReady;
  assign execute_ctrl10_down_LANE_SEL_lane0 = execute_ctrl10_up_LANE_SEL_lane0;
  assign execute_ctrl10_down_TRAP_lane0 = execute_ctrl10_up_TRAP_lane0;
  assign execute_ctrl10_down_Decode_UOP_ID_lane0 = execute_ctrl10_up_Decode_UOP_ID_lane0;
  assign execute_ctrl10_down_RD_ENABLE_lane0 = execute_ctrl10_up_RD_ENABLE_lane0;
  assign execute_ctrl10_down_RD_RFID_lane0 = execute_ctrl10_up_RD_RFID_lane0;
  assign execute_ctrl10_down_RD_PHYS_lane0 = execute_ctrl10_up_RD_PHYS_lane0;
  assign execute_ctrl10_down_LANE_AGE_lane0 = execute_ctrl10_up_LANE_AGE_lane0;
  assign execute_ctrl10_down_COMPLETED_lane0 = execute_ctrl10_up_COMPLETED_lane0;
  assign execute_ctrl10_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl10_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl10_down_COMPLETION_AT_11_lane0 = execute_ctrl10_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl10_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl10_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl10_down_COMMIT_lane0 = execute_ctrl10_up_COMMIT_lane0;
  assign execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl10_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  assign execute_ctrl11_up_ready = execute_ctrl11_down_isReady;
  assign execute_ctrl11_down_LANE_SEL_lane0 = execute_ctrl11_up_LANE_SEL_lane0;
  assign execute_ctrl11_down_TRAP_lane0 = execute_ctrl11_up_TRAP_lane0;
  assign execute_ctrl11_down_Decode_UOP_ID_lane0 = execute_ctrl11_up_Decode_UOP_ID_lane0;
  assign execute_ctrl11_down_RD_ENABLE_lane0 = execute_ctrl11_up_RD_ENABLE_lane0;
  assign execute_ctrl11_down_RD_RFID_lane0 = execute_ctrl11_up_RD_RFID_lane0;
  assign execute_ctrl11_down_RD_PHYS_lane0 = execute_ctrl11_up_RD_PHYS_lane0;
  assign execute_ctrl11_down_LANE_AGE_lane0 = execute_ctrl11_up_LANE_AGE_lane0;
  assign execute_ctrl11_down_lane0_float_WriteBackPlugin_SEL_lane0 = execute_ctrl11_up_lane0_float_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl11_down_COMPLETION_AT_11_lane0 = execute_ctrl11_up_COMPLETION_AT_11_lane0;
  assign execute_ctrl11_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl11_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl11_down_COMMIT_lane0 = execute_ctrl11_up_COMMIT_lane0;
  assign execute_ctrl12_up_ready = execute_ctrl12_down_isReady;
  assign execute_ctrl12_down_RD_RFID_lane0 = execute_ctrl12_up_RD_RFID_lane0;
  assign execute_ctrl12_down_RD_PHYS_lane0 = execute_ctrl12_up_RD_PHYS_lane0;
  assign execute_ctrl12_down_LANE_AGE_lane0 = execute_ctrl12_up_LANE_AGE_lane0;
  assign execute_ctrl12_down_lane0_float_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl12_up_lane0_float_WriteBackPlugin_logic_DATA_lane0;
  assign fetch_logic_ctrls_0_down_isFiring = (fetch_logic_ctrls_0_down_isValid && fetch_logic_ctrls_0_down_isReady);
  assign fetch_logic_ctrls_0_down_isValid = fetch_logic_ctrls_0_down_valid;
  assign fetch_logic_ctrls_0_down_isReady = fetch_logic_ctrls_0_down_ready;
  assign fetch_logic_ctrls_1_up_isValid = fetch_logic_ctrls_1_up_valid;
  assign fetch_logic_ctrls_1_up_isReady = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_up_isCancel = fetch_logic_ctrls_1_up_cancel;
  assign fetch_logic_ctrls_1_down_isValid = fetch_logic_ctrls_1_down_valid;
  assign fetch_logic_ctrls_1_down_isReady = fetch_logic_ctrls_1_down_ready;
  assign fetch_logic_ctrls_2_up_isValid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_isReady = fetch_logic_ctrls_2_up_ready;
  assign fetch_logic_ctrls_2_up_isCancel = fetch_logic_ctrls_2_up_cancel;
  assign fetch_logic_ctrls_2_up_isCanceling = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isCancel);
  assign fetch_logic_ctrls_0_up_isFiring = (fetch_logic_ctrls_0_up_isValid && fetch_logic_ctrls_0_up_isReady);
  assign fetch_logic_ctrls_0_up_isValid = fetch_logic_ctrls_0_up_valid;
  assign fetch_logic_ctrls_0_up_isReady = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_2_down_isValid = fetch_logic_ctrls_2_down_valid;
  assign fetch_logic_ctrls_2_down_isReady = fetch_logic_ctrls_2_down_ready;
  assign fetch_logic_ctrls_2_down_isCancel = 1'b0;
  assign decode_ctrls_0_down_isValid = decode_ctrls_0_down_valid;
  assign decode_ctrls_0_down_isReady = decode_ctrls_0_down_ready;
  assign decode_ctrls_1_up_isMoving = (decode_ctrls_1_up_isValid && decode_ctrls_1_up_isReady);
  assign decode_ctrls_1_up_isValid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_isReady = decode_ctrls_1_up_ready;
  assign decode_ctrls_1_up_isCanceling = 1'b0;
  assign decode_ctrls_0_up_isFiring = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isMoving = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isValid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_isReady = decode_ctrls_0_up_ready;
  assign decode_ctrls_0_up_isCancel = 1'b0;
  assign decode_ctrls_1_down_isReady = decode_ctrls_1_down_ready;
  assign execute_ctrl0_down_isReady = execute_ctrl0_down_ready;
  assign execute_ctrl1_down_isReady = execute_ctrl1_down_ready;
  assign execute_ctrl2_down_isReady = execute_ctrl2_down_ready;
  assign execute_ctrl3_down_isReady = execute_ctrl3_down_ready;
  assign execute_ctrl4_down_isReady = execute_ctrl4_down_ready;
  assign execute_ctrl5_down_isReady = execute_ctrl5_down_ready;
  assign execute_ctrl6_down_isReady = execute_ctrl6_down_ready;
  assign execute_ctrl7_down_isReady = execute_ctrl7_down_ready;
  assign execute_ctrl8_down_isReady = execute_ctrl8_down_ready;
  assign execute_ctrl9_down_isReady = execute_ctrl9_down_ready;
  assign execute_ctrl10_down_isReady = execute_ctrl10_down_ready;
  assign execute_ctrl11_down_isReady = execute_ctrl11_down_ready;
  assign execute_ctrl12_down_isReady = execute_ctrl12_down_ready;
  always @(*) begin
    LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_stateReg;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_SB_DRAIN : begin
        if(LsuPlugin_logic_storeBuffer_empty) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_CMD;
        end
      end
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l363) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_COMPLETION;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l371) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
        end
      end
      default : begin
        if(LsuPlugin_logic_flusher_arbiter_io_output_valid) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_SB_DRAIN;
        end
      end
    endcase
    if(LsuPlugin_logic_flusher_wantKill) begin
      LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
    end
  end

  assign when_LsuPlugin_l363 = (LsuPlugin_logic_flusher_cmdCounter[6] && (! LsuPlugin_logic_flusher_inflight));
  assign when_LsuPlugin_l371 = (! (|LsuPlugin_logic_flusher_waiter));
  assign LsuPlugin_logic_flusher_onExit_IDLE = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onExit_SB_DRAIN = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_SB_DRAIN) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_SB_DRAIN));
  assign LsuPlugin_logic_flusher_onExit_CMD = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onExit_COMPLETION = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_COMPLETION));
  assign LsuPlugin_logic_flusher_onEntry_IDLE = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onEntry_SB_DRAIN = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_SB_DRAIN) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_SB_DRAIN));
  assign LsuPlugin_logic_flusher_onEntry_CMD = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onEntry_COMPLETION = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_COMPLETION));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_stateReg;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_COMPUTE;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        if(when_TrapPlugin_l409) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL;
        end else begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
            end
            4'b0001 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC;
            end
            4'b0010 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH;
            end
            4'b0100 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b0101 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b1000 : begin
              if(TrapPlugin_api_harts_0_askWake) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
              end
            end
            4'b0110 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        if(TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        if(TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
        end
      end
      default : begin
        if(when_TrapPlugin_l362) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
        end
      end
    endcase
    if(TrapPlugin_logic_harts_0_trap_fsm_wantKill) begin
      TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RESET;
    end
  end

  assign when_TrapPlugin_l409 = ((TrapPlugin_logic_harts_0_trap_pending_state_exception || TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak) || TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt);
  assign when_TrapPlugin_l654 = (TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege != 2'b11);
  assign switch_TrapPlugin_l655 = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign when_TrapPlugin_l362 = (&TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0);
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_COMPUTE = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_COMPUTE) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_COMPUTE));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_COMPUTE = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_COMPUTE) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_COMPUTE));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  always @(*) begin
    CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_stateReg;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l296) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_WRITE;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l325) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_COMPLETION;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
        end
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(when_CsrAccessPlugin_l212) begin
            CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
          end
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
            end
          end
        end
      end
    endcase
    if(CsrAccessPlugin_logic_fsm_wantKill) begin
      CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
    end
  end

  assign when_CsrAccessPlugin_l296 = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l325 = (! CsrAccessPlugin_bus_write_halt);
  assign when_CsrAccessPlugin_l212 = ((! CsrAccessPlugin_logic_fsm_inject_trap) && (! CsrAccessPlugin_bus_decode_trap));
  assign CsrAccessPlugin_logic_fsm_onExit_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onExit_READ = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onExit_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onExit_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_COMPLETION));
  assign CsrAccessPlugin_logic_fsm_onEntry_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onEntry_READ = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onEntry_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onEntry_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_COMPLETION));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      FpuCsrPlugin_api_rm <= 3'b000;
      LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      LsuL1Plugin_logic_refill_slots_1_valid <= 1'b0;
      LsuL1Plugin_logic_refill_slots_1_loaded <= 1'b1;
      LsuL1Plugin_logic_refill_pushCounter <= 32'h0;
      LsuL1Plugin_logic_refill_read_arbiter_lock <= 2'b00;
      LsuL1Plugin_logic_refill_read_wordIndex <= 1'b0;
      LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_busy <= 1'b0;
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= 2'b00;
      LsuL1Plugin_logic_writeback_read_wordIndex <= 1'b0;
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= 2'b00;
      LsuL1Plugin_logic_writeback_write_wordIndex <= 1'b0;
      LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= 1'b0;
      LsuL1Plugin_logic_initializer_counter <= 7'h0;
      PrefetcherRptPlugin_logic_csr_disable <= 1'b0;
      PrefetcherRptPlugin_logic_counter <= 3'b000;
      PrefetcherRptPlugin_logic_pip2_node_1_valid <= 1'b0;
      _zz_25 <= 1'b0;
      PrivilegedPlugin_logic_harts_0_privilege <= 2'b11;
      PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_fs <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_meie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_mtie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_msie <= 1'b0;
      FpuCsrPlugin_api_flags_NV <= 1'b0;
      FpuCsrPlugin_api_flags_DZ <= 1'b0;
      FpuCsrPlugin_api_flags_OF <= 1'b0;
      FpuCsrPlugin_api_flags_UF <= 1'b0;
      FpuCsrPlugin_api_flags_NX <= 1'b0;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_counter <= 1'b0;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rValid <= 1'b0;
      FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      FetchL1Plugin_logic_invalidate_firstEver <= 1'b1;
      FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      FetchL1Plugin_logic_refill_slots_1_valid <= 1'b0;
      FetchL1Plugin_logic_refill_slots_1_cmdSent <= 1'b1;
      FetchL1Plugin_logic_refill_pushCounter <= 32'h0;
      FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      FetchL1Plugin_logic_refill_onRsp_wordIndex <= 1'b0;
      FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= 1'b0;
      FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      BtbPlugin_logic_ras_ptr_push <= 2'b00;
      BtbPlugin_logic_ras_ptr_pop <= 2'b11;
      decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      decode_ctrls_0_up_LANE_SEL_1_regNext <= 1'b0;
      FetchL1Plugin_logic_bus_toWishbone_counter <= 1'b0;
      _zz_FetchL1Plugin_logic_bus_rsp_valid <= 1'b0;
      FpuAddSharedPlugin_logic_pip_node_1_valid <= 1'b0;
      FpuAddSharedPlugin_logic_pip_node_2_valid <= 1'b0;
      FpuAddSharedPlugin_logic_pip_node_3_valid <= 1'b0;
      FpuAddSharedPlugin_logic_pip_node_4_valid <= 1'b0;
      early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      AlignerPlugin_logic_feeder_harts_0_dopId <= 10'h0;
      AlignerPlugin_logic_buffer_mask <= 4'b0000;
      AlignerPlugin_logic_buffer_last <= 4'b0000;
      AlignerPlugin_logic_buffer_trap <= 1'b0;
      LsuPlugin_logic_storeBuffer_ops_pushPtr <= 6'h0;
      LsuPlugin_logic_storeBuffer_ops_popPtr <= 6'h0;
      LsuPlugin_logic_storeBuffer_ops_freePtr <= 6'h0;
      LsuPlugin_logic_storeBuffer_slots_0_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_1_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_2_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_3_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_4_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_5_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_6_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_slots_7_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_holdHart_waitIt <= 1'b0;
      LsuPlugin_logic_storeBuffer_waitL1_valid <= 1'b0;
      LsuPlugin_logic_onAddress0_ls_storeId <= 12'h0;
      execute_ctrl3_up_LsuL1_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LsuL1_SEL_lane0 <= 1'b0;
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      LsuPlugin_logic_onCtrl_io_doItReg <= 1'b0;
      LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      LsuPlugin_logic_onCtrl_commitProbeToken <= 1'b0;
      LsuPlugin_logic_storeBuffer_ops_pip_node_1_valid <= 1'b0;
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_valid <= 1'b0;
      FpuPackerPlugin_logic_s1_subnormal_counter <= 2'b00;
      FpuPackerPlugin_logic_pip_node_1_valid <= 1'b0;
      FpuPackerPlugin_logic_pip_node_2_valid <= 1'b0;
      LsuPlugin_logic_bus_cmd_rValid <= 1'b0;
      PrefetcherRptPlugin_logic_pip_node_1_valid <= 1'b0;
      PrefetcherRptPlugin_logic_pip_node_2_valid <= 1'b0;
      CsrRamPlugin_csrMapper_fired <= 1'b0;
      late0_BranchPlugin_logic_jumpLogic_learn_rValid <= 1'b0;
      late1_BranchPlugin_logic_jumpLogic_learn_rValid <= 1'b0;
      DecoderPlugin_logic_harts_0_uopId <= 16'h0;
      DecoderPlugin_logic_interrupt_buffered <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_1_regNext <= 1'b0;
      DispatchPlugin_logic_slots_0_ctx_valid <= 1'b0;
      DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      DispatchPlugin_logic_feeds_1_sent <= 1'b0;
      FpuUnpack_RS1_normalizer_validReg <= 1'b0;
      FpuUnpack_RS1_normalizer_asked <= 1'b0;
      FpuUnpack_RS1_normalizer_served <= 1'b0;
      FpuUnpack_RS2_normalizer_validReg <= 1'b0;
      FpuUnpack_RS2_normalizer_asked <= 1'b0;
      FpuUnpack_RS2_normalizer_served <= 1'b0;
      FpuUnpack_RS3_normalizer_validReg <= 1'b0;
      FpuUnpack_RS3_normalizer_asked <= 1'b0;
      FpuUnpack_RS3_normalizer_served <= 1'b0;
      FpuUnpackerPlugin_logic_onCvt_asked <= 1'b0;
      FpuUnpackerPlugin_logic_onCvt_served <= 1'b0;
      FpuUnpackerPlugin_logic_unpacker_node_1_valid <= 1'b0;
      FpuUnpackerPlugin_logic_unpacker_node_2_valid <= 1'b0;
      FpuF2iPlugin_logic_onResult_halfRater_firstCycle <= 1'b1;
      FpuSqrtPlugin_logic_onExecute_isZero <= 1'b0;
      FpuSqrtPlugin_logic_onExecute_cmdSent <= 1'b0;
      FpuSqrtPlugin_logic_onExecute_unscheduleRequest <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= 1'b0;
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      execute_ctrl0_down_LANE_SEL_lane1_regNext <= 1'b0;
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      execute_ctrl2_down_LANE_SEL_lane1_regNext <= 1'b0;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_1 <= 1'b0;
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
      PcPlugin_logic_harts_0_self_id <= 10'h0;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      PcPlugin_logic_harts_0_self_fault <= 1'b0;
      PcPlugin_logic_harts_0_self_state <= 32'h0;
      PcPlugin_logic_harts_0_holdReg <= 1'b1;
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_sampled <= 1'b0;
      HistoryPlugin_logic_onFetch_value <= 12'h0;
      CsrRamPlugin_logic_readLogic_ohReg <= 2'b00;
      CsrRamPlugin_logic_readLogic_busy <= 1'b0;
      CsrRamPlugin_logic_flush_counter <= 3'b000;
      execute_ctrl1_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl2_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl3_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl5_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl6_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl7_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl8_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl9_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl10_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl11_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl12_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl1_up_LANE_SEL_lane1 <= 1'b0;
      execute_ctrl2_up_LANE_SEL_lane1 <= 1'b0;
      execute_ctrl3_up_LANE_SEL_lane1 <= 1'b0;
      execute_ctrl4_up_LANE_SEL_lane1 <= 1'b0;
      execute_ctrl5_up_LANE_SEL_lane1 <= 1'b0;
      integer_RegFilePlugin_logic_initalizer_counter <= 6'h0;
      float_RegFilePlugin_logic_initalizer_counter <= 6'h0;
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 <= 60'h0;
      fetch_logic_ctrls_1_up_valid <= 1'b0;
      fetch_logic_ctrls_2_up_valid <= 1'b0;
      decode_ctrls_1_up_valid <= 1'b0;
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_IDLE;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_RESET;
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_IDLE;
    end else begin
      if(LsuL1Plugin_logic_refill_slots_0_loadedSet) begin
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_0_fire) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_refill_slots_1_loadedSet) begin
        LsuL1Plugin_logic_refill_slots_1_loaded <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_1_fire) begin
        LsuL1Plugin_logic_refill_slots_1_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_refill_push_valid) begin
        LsuL1Plugin_logic_refill_pushCounter <= (LsuL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(when_LsuL1Plugin_l377) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b0;
      end
      if(when_LsuL1Plugin_l377_1) begin
        LsuL1Plugin_logic_refill_slots_1_valid <= 1'b1;
        LsuL1Plugin_logic_refill_slots_1_loaded <= 1'b0;
      end
      LsuL1Plugin_logic_refill_read_arbiter_lock <= LsuL1Plugin_logic_refill_read_arbiter_oh;
      if(LsuL1Plugin_logic_bus_read_cmd_fire) begin
        LsuL1Plugin_logic_refill_read_arbiter_lock <= 2'b00;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_writeReservation_win); // LsuL1Plugin.scala:L429
          `else
            if(!LsuL1Plugin_logic_refill_read_writeReservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L429
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l450) begin
        LsuL1Plugin_logic_refill_read_hadError <= 1'b1;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_reservation_win); // LsuL1Plugin.scala:L459
          `else
            if(!LsuL1Plugin_logic_refill_read_reservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L459
              $finish;
            end
          `endif
        `endif
        if(LsuL1Plugin_logic_refill_read_rspWithData) begin
          LsuL1Plugin_logic_refill_read_wordIndex <= (LsuL1Plugin_logic_refill_read_wordIndex + 1'b1);
        end
        if(when_LsuL1Plugin_l463) begin
          LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
        end
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      end
      if(when_LsuL1Plugin_l530) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_slots_1_fire) begin
        LsuL1Plugin_logic_writeback_slots_1_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_slots_1_fire) begin
        LsuL1Plugin_logic_writeback_slots_1_busy <= 1'b0;
      end
      if(when_LsuL1Plugin_l530_1) begin
        LsuL1Plugin_logic_writeback_slots_1_valid <= 1'b0;
      end
      if(when_LsuL1Plugin_l556) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b1;
      end
      if(when_LsuL1Plugin_l556_1) begin
        LsuL1Plugin_logic_writeback_slots_1_valid <= 1'b1;
        LsuL1Plugin_logic_writeback_slots_1_busy <= 1'b1;
      end
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= LsuL1Plugin_logic_writeback_read_arbiter_oh;
      LsuL1Plugin_logic_writeback_read_wordIndex <= (LsuL1Plugin_logic_writeback_read_wordIndex + LsuL1Plugin_logic_writeback_read_slotRead_valid);
      if(when_LsuL1Plugin_l605) begin
        LsuL1Plugin_logic_writeback_read_arbiter_lock <= 2'b00;
      end
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= LsuL1Plugin_logic_writeback_read_slotRead_valid;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= LsuL1Plugin_logic_writeback_write_arbiter_oh;
      LsuL1Plugin_logic_writeback_write_wordIndex <= (LsuL1Plugin_logic_writeback_write_wordIndex + (LsuL1Plugin_logic_writeback_write_bufferRead_fire && 1'b1));
      if(when_LsuL1Plugin_l676) begin
        LsuL1Plugin_logic_writeback_write_arbiter_lock <= 2'b00;
      end
      if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
        LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= LsuL1Plugin_logic_writeback_write_bufferRead_valid;
      end
      if(LsuL1Plugin_logic_banks_0_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_1_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735_1) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      end
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= (execute_ctrl4_down_LsuL1_HAZARD_lane0 && execute_freeze_valid);
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= (execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 && execute_freeze_valid);
      if(execute_ctrl4_down_LsuL1_SEL_lane0) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_59 <= 2'b01)); // LsuL1Plugin.scala:L892
          `else
            if(!(_zz_59 <= 2'b01)) begin
              $display("FAILURE Multiple way hit ???"); // LsuL1Plugin.scala:L892
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l915) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_61 < 2'b10)); // LsuL1Plugin.scala:L916
          `else
            if(!(_zz_61 < 2'b10)) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L916
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l1218) begin
        LsuL1Plugin_logic_initializer_counter <= (LsuL1Plugin_logic_initializer_counter + 7'h01);
      end
      PrefetcherRptPlugin_logic_counter <= ((! PrefetcherRptPlugin_logic_queued_ready) ? _zz_PrefetcherRptPlugin_logic_counter : 3'b000);
      if(PrefetcherRptPlugin_logic_pip2_node_0_isReady) begin
        PrefetcherRptPlugin_logic_pip2_node_1_valid <= PrefetcherRptPlugin_logic_pip2_node_0_isValid;
      end
      _zz_25 <= (! PrefetcherRptPlugin_logic_order_ready);
      if(PrivilegedPlugin_logic_harts_0_xretAwayFromMachine) begin
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      end
      if(when_PrivilegedPlugin_l550) begin
        PrivilegedPlugin_logic_harts_0_m_status_fs <= 2'b11;
      end
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= PrivilegedPlugin_logic_harts_0_int_m_external;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= PrivilegedPlugin_logic_harts_0_int_m_timer;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= PrivilegedPlugin_logic_harts_0_int_m_software;
      if(LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_fire) begin
        LsuL1Plugin_logic_bus_toWishbone_arbiter_counter <= (LsuL1Plugin_logic_bus_toWishbone_arbiter_counter + 1'b1);
      end
      if(LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready) begin
        LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rValid <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_valid;
      end
      if(FetchL1Plugin_logic_invalidate_done) begin
        FetchL1Plugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchL1Plugin_l204) begin
        FetchL1Plugin_logic_invalidate_counter <= FetchL1Plugin_logic_invalidate_counterIncr;
      end
      if(when_FetchL1Plugin_l211) begin
        FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      end
      if(when_FetchL1Plugin_l255) begin
        if(_zz_38) begin
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
        end
        if(_zz_when) begin
          FetchL1Plugin_logic_refill_slots_1_valid <= 1'b1;
          FetchL1Plugin_logic_refill_slots_1_cmdSent <= 1'b0;
        end
        FetchL1Plugin_logic_refill_pushCounter <= (FetchL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(FetchL1Plugin_logic_bus_cmd_valid) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b1;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        if(_zz_FetchL1Plugin_logic_bus_cmd_payload_address) begin
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
        end
        if(_zz_FetchL1Plugin_logic_bus_cmd_payload_id) begin
          FetchL1Plugin_logic_refill_slots_1_cmdSent <= 1'b1;
        end
      end
      if(FetchL1Plugin_logic_bus_rsp_fire) begin
        FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_rsp_valid) begin
        FetchL1Plugin_logic_refill_onRsp_wordIndex <= (FetchL1Plugin_logic_refill_onRsp_wordIndex + 1'b1);
        if(when_FetchL1Plugin_l330) begin
          FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
          case(FetchL1Plugin_logic_bus_rsp_payload_id)
            1'b0 : begin
              FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
            end
            default : begin
              FetchL1Plugin_logic_refill_slots_1_valid <= 1'b0;
            end
          endcase
        end
      end
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
      if(FetchL1Plugin_logic_trapPort_valid) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b1;
      end
      if(fetch_logic_ctrls_2_up_isCancel) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      end
      if(fetch_logic_ctrls_2_up_isValid) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b0;
      end
      if(when_FetchL1Plugin_l541) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((|{FetchL1Plugin_logic_refill_slots_1_valid,FetchL1Plugin_logic_refill_slots_0_valid}) && (! FetchL1Plugin_logic_invalidate_done)))); // FetchL1Plugin.scala:L556
        `else
          if(!(! ((|{FetchL1Plugin_logic_refill_slots_1_valid,FetchL1Plugin_logic_refill_slots_0_valid}) && (! FetchL1Plugin_logic_invalidate_done)))) begin
            $display("FAILURE "); // FetchL1Plugin.scala:L556
            $finish;
          end
        `endif
      `endif
      BtbPlugin_logic_ras_ptr_push <= (_zz_BtbPlugin_logic_ras_ptr_push - _zz_BtbPlugin_logic_ras_ptr_push_3);
      decode_ctrls_0_up_LANE_SEL_0_regNext <= decode_ctrls_0_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50) begin
        decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      end
      decode_ctrls_0_up_LANE_SEL_1_regNext <= decode_ctrls_0_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l50_1) begin
        decode_ctrls_0_up_LANE_SEL_1_regNext <= 1'b0;
      end
      if(when_FetchL1Bus_l247) begin
        if(when_FetchL1Bus_l250) begin
          FetchL1Plugin_logic_bus_toWishbone_counter <= (FetchL1Plugin_logic_bus_toWishbone_counter + 1'b1);
        end
      end
      _zz_FetchL1Plugin_logic_bus_rsp_valid <= (FetchL1WishbonePlugin_logic_bus_CYC && (FetchL1WishbonePlugin_logic_bus_ACK || FetchL1WishbonePlugin_logic_bus_ERR));
      if(FpuAddSharedPlugin_logic_pip_node_0_isValid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_63 <= 2'b01)); // FpuAddSharedPlugin.scala:L108
          `else
            if(!(_zz_63 <= 2'b01)) begin
              $display("FAILURE "); // FpuAddSharedPlugin.scala:L108
              $finish;
            end
          `endif
        `endif
      end
      if(FpuAddSharedPlugin_logic_pip_node_0_isReady) begin
        FpuAddSharedPlugin_logic_pip_node_1_valid <= FpuAddSharedPlugin_logic_pip_node_0_isValid;
      end
      if(FpuAddSharedPlugin_logic_pip_node_1_isReady) begin
        FpuAddSharedPlugin_logic_pip_node_2_valid <= FpuAddSharedPlugin_logic_pip_node_1_isValid;
      end
      if(FpuAddSharedPlugin_logic_pip_node_2_isReady) begin
        FpuAddSharedPlugin_logic_pip_node_3_valid <= FpuAddSharedPlugin_logic_pip_node_2_isValid;
      end
      if(FpuAddSharedPlugin_logic_pip_node_3_isReady) begin
        FpuAddSharedPlugin_logic_pip_node_4_valid <= FpuAddSharedPlugin_logic_pip_node_3_isValid;
      end
      if(io_cmd_fire) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      end
      early0_DivPlugin_logic_processing_unscheduleRequest <= execute_lane0_ctrls_2_upIsCancel;
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      end
      if(when_AlignerPlugin_l171) begin
        AlignerPlugin_logic_feeder_harts_0_dopId <= (decode_ctrls_0_down_Decode_DOP_ID_1 + 10'h001);
      end
      if(AlignerPlugin_logic_buffer_downFire) begin
        AlignerPlugin_logic_buffer_mask <= (AlignerPlugin_logic_buffer_mask & (~ AlignerPlugin_logic_buffer_usedMask[3 : 0]));
        AlignerPlugin_logic_buffer_last <= (AlignerPlugin_logic_buffer_last & (~ AlignerPlugin_logic_buffer_usedMask[3 : 0]));
      end
      if(when_AlignerPlugin_l256) begin
        AlignerPlugin_logic_buffer_mask <= (fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[7 : 4] : 4'b0000)));
        AlignerPlugin_logic_buffer_trap <= fetch_logic_ctrls_2_down_TRAP;
        AlignerPlugin_logic_buffer_last <= fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
      end
      LsuPlugin_logic_storeBuffer_ops_popPtr <= (LsuPlugin_logic_storeBuffer_ops_popPtr + _zz_LsuPlugin_logic_storeBuffer_ops_popPtr);
      if(LsuPlugin_logic_storeBuffer_push_valid) begin
        LsuPlugin_logic_storeBuffer_ops_pushPtr <= (LsuPlugin_logic_storeBuffer_ops_pushPtr + _zz_LsuPlugin_logic_storeBuffer_ops_pushPtr);
        if(_zz_when_3) begin
          LsuPlugin_logic_storeBuffer_slots_0_valid <= 1'b1;
        end
        if(_zz_when_4) begin
          LsuPlugin_logic_storeBuffer_slots_1_valid <= 1'b1;
        end
        if(_zz_when_5) begin
          LsuPlugin_logic_storeBuffer_slots_2_valid <= 1'b1;
        end
        if(_zz_when_6) begin
          LsuPlugin_logic_storeBuffer_slots_3_valid <= 1'b1;
        end
        if(_zz_when_7) begin
          LsuPlugin_logic_storeBuffer_slots_4_valid <= 1'b1;
        end
        if(_zz_when_8) begin
          LsuPlugin_logic_storeBuffer_slots_5_valid <= 1'b1;
        end
        if(_zz_when_9) begin
          LsuPlugin_logic_storeBuffer_slots_6_valid <= 1'b1;
        end
        if(_zz_when_10) begin
          LsuPlugin_logic_storeBuffer_slots_7_valid <= 1'b1;
        end
      end
      if(when_LsuPlugin_l331) begin
        LsuPlugin_logic_storeBuffer_holdHart_waitIt <= 1'b0;
      end
      if(when_LsuPlugin_l259) begin
        LsuPlugin_logic_storeBuffer_waitL1_valid <= 1'b0;
      end
      LsuPlugin_logic_onAddress0_ls_storeId <= (LsuPlugin_logic_onAddress0_ls_storeId + _zz_LsuPlugin_logic_onAddress0_ls_storeId);
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b1;
      if(execute_freeze_valid) begin
        LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      if(when_LsuPlugin_l597) begin
        LsuPlugin_logic_onCtrl_io_allowIt <= 1'b1;
      end
      LsuPlugin_logic_onCtrl_io_doItReg <= LsuPlugin_logic_onCtrl_io_doIt;
      if(LsuPlugin_logic_bus_cmd_fire) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b1;
      end
      if(when_LsuPlugin_l601) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      end
      if(LsuPlugin_logic_bus_rsp_toStream_valid) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b1;
      end
      if(LsuPlugin_logic_onCtrl_io_rsp_fire) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      end
      if(when_LsuPlugin_l686) begin
        if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
        end
      end
      if(when_LsuPlugin_l705) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      end
      if(when_LsuPlugin_l709) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
      end
      if(when_LsuPlugin_l865) begin
        if(when_LsuPlugin_l876) begin
          LsuPlugin_logic_storeBuffer_holdHart_waitIt <= 1'b1;
        end
      end
      if(when_LsuPlugin_l910) begin
        if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
          LsuPlugin_logic_storeBuffer_ops_popPtr <= LsuPlugin_logic_storeBuffer_ops_freePtr;
          if(when_LsuPlugin_l913) begin
            if(when_LsuPlugin_l263) begin
              LsuPlugin_logic_storeBuffer_waitL1_valid <= 1'b1;
            end
          end
        end else begin
          LsuPlugin_logic_storeBuffer_ops_freePtr <= (LsuPlugin_logic_storeBuffer_ops_freePtr + 6'h01);
          if(when_LsuPlugin_l918) begin
            LsuPlugin_logic_storeBuffer_slots_0_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_1) begin
            LsuPlugin_logic_storeBuffer_slots_1_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_2) begin
            LsuPlugin_logic_storeBuffer_slots_2_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_3) begin
            LsuPlugin_logic_storeBuffer_slots_3_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_4) begin
            LsuPlugin_logic_storeBuffer_slots_4_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_5) begin
            LsuPlugin_logic_storeBuffer_slots_5_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_6) begin
            LsuPlugin_logic_storeBuffer_slots_6_valid <= 1'b0;
          end
          if(when_LsuPlugin_l918_7) begin
            LsuPlugin_logic_storeBuffer_slots_7_valid <= 1'b0;
          end
        end
      end
      if(when_LsuPlugin_l259_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      end
      if(when_LsuPlugin_l949) begin
        if(when_LsuPlugin_l263_1) begin
          LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b1;
        end
      end
      if(LsuPlugin_logic_onCtrl_commitProbeReq) begin
        LsuPlugin_logic_onCtrl_commitProbeToken <= LsuPlugin_logic_onCtrl_lsuTrap;
      end
      if(LsuPlugin_logic_storeBuffer_ops_pip_node_0_isReady) begin
        LsuPlugin_logic_storeBuffer_ops_pip_node_1_valid <= LsuPlugin_logic_storeBuffer_ops_pip_node_0_isValid;
      end
      if(LsuPlugin_logic_storeBuffer_ops_pip_node_1_isReady) begin
        LsuPlugin_logic_storeBuffer_ops_pip_node_2_valid <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_isValid;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((_zz_65 <= 3'b001)); // FpuPackerPlugin.scala:L104
        `else
          if(!(_zz_65 <= 3'b001)) begin
            $display("FAILURE Packing GROUP_OH failure"); // FpuPackerPlugin.scala:L104
            $finish;
          end
        `endif
      `endif
      if(FpuPackerPlugin_logic_s1_subnormal_freezeIt) begin
        FpuPackerPlugin_logic_s1_subnormal_counter <= (FpuPackerPlugin_logic_s1_subnormal_counter + 2'b01);
      end
      if(when_FpuPackerPlugin_l134) begin
        FpuPackerPlugin_logic_s1_subnormal_counter <= 2'b00;
      end
      if(FpuPackerPlugin_logic_pip_node_0_isReady) begin
        FpuPackerPlugin_logic_pip_node_1_valid <= FpuPackerPlugin_logic_pip_node_0_isValid;
      end
      if(FpuPackerPlugin_logic_pip_node_1_isReady) begin
        FpuPackerPlugin_logic_pip_node_2_valid <= FpuPackerPlugin_logic_pip_node_1_isValid;
      end
      if(LsuPlugin_logic_bus_cmd_ready) begin
        LsuPlugin_logic_bus_cmd_rValid <= LsuPlugin_logic_bus_cmd_valid;
      end
      PrefetcherRptPlugin_logic_pip_node_1_valid <= PrefetcherRptPlugin_logic_pip_node_0_isValid;
      PrefetcherRptPlugin_logic_pip_node_2_valid <= PrefetcherRptPlugin_logic_pip_node_1_isValid;
      if(when_CsrRamPlugin_l92) begin
        CsrRamPlugin_csrMapper_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        CsrRamPlugin_csrMapper_fired <= 1'b0;
      end
      if(late0_BranchPlugin_logic_jumpLogic_learn_ready) begin
        late0_BranchPlugin_logic_jumpLogic_learn_rValid <= late0_BranchPlugin_logic_jumpLogic_learn_valid;
      end
      if(late1_BranchPlugin_logic_jumpLogic_learn_ready) begin
        late1_BranchPlugin_logic_jumpLogic_learn_rValid <= late1_BranchPlugin_logic_jumpLogic_learn_valid;
      end
      if(when_DecoderPlugin_l143) begin
        DecoderPlugin_logic_harts_0_uopId <= (DecoderPlugin_logic_harts_0_uopId + 16'h0002);
      end
      if(when_DecoderPlugin_l151) begin
        DecoderPlugin_logic_interrupt_buffered <= DecoderPlugin_logic_interrupt_async;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_2) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      end
      decode_ctrls_1_up_LANE_SEL_1_regNext <= decode_ctrls_1_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l50_3) begin
        decode_ctrls_1_up_LANE_SEL_1_regNext <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_0_sending) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b1;
      end
      if(decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_1_sending) begin
        DispatchPlugin_logic_feeds_1_sent <= 1'b1;
      end
      if(decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_1_sent <= 1'b0;
      end
      if(when_DispatchPlugin_l378) begin
        DispatchPlugin_logic_slots_0_ctx_valid <= 1'b0;
      end
      FpuUnpack_RS1_normalizer_validReg <= (FpuUnpack_RS1_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0);
      if(when_FpuUnpackerPlugin_l234) begin
        FpuUnpack_RS1_normalizer_validReg <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l235) begin
        FpuUnpack_RS1_normalizer_asked <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS1_normalizer_asked <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l236) begin
        FpuUnpack_RS1_normalizer_served <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS1_normalizer_served <= 1'b0;
      end
      FpuUnpack_RS2_normalizer_validReg <= (FpuUnpack_RS2_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS2_IS_SUBNORMAL_lane0);
      if(when_FpuUnpackerPlugin_l234_1) begin
        FpuUnpack_RS2_normalizer_validReg <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l235_1) begin
        FpuUnpack_RS2_normalizer_asked <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS2_normalizer_asked <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l236_1) begin
        FpuUnpack_RS2_normalizer_served <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS2_normalizer_served <= 1'b0;
      end
      FpuUnpack_RS3_normalizer_validReg <= (FpuUnpack_RS3_normalizer_unpackerSel && execute_ctrl2_down_FpuUnpack_RS3_IS_SUBNORMAL_lane0);
      if(when_FpuUnpackerPlugin_l234_2) begin
        FpuUnpack_RS3_normalizer_validReg <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l235_2) begin
        FpuUnpack_RS3_normalizer_asked <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS3_normalizer_asked <= 1'b0;
      end
      if(when_FpuUnpackerPlugin_l236_2) begin
        FpuUnpack_RS3_normalizer_served <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpack_RS3_normalizer_served <= 1'b0;
      end
      if(FpuUnpackerPlugin_logic_unpacker_arbiter_io_inputs_1_ready) begin
        FpuUnpackerPlugin_logic_onCvt_asked <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpackerPlugin_logic_onCvt_asked <= 1'b0;
      end
      if(FpuUnpackerPlugin_logic_unpacker_results_1_valid) begin
        FpuUnpackerPlugin_logic_onCvt_served <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuUnpackerPlugin_logic_onCvt_served <= 1'b0;
      end
      FpuUnpackerPlugin_logic_unpacker_node_1_valid <= FpuUnpackerPlugin_logic_unpacker_node_0_isValid;
      FpuUnpackerPlugin_logic_unpacker_node_2_valid <= FpuUnpackerPlugin_logic_unpacker_node_1_isValid;
      FpuF2iPlugin_logic_onResult_halfRater_firstCycle <= (! execute_freeze_valid);
      if(when_FpuSqrtPlugin_l66) begin
        FpuSqrtPlugin_logic_onExecute_isZero <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuSqrtPlugin_logic_onExecute_isZero <= 1'b0;
      end
      if(io_input_fire) begin
        FpuSqrtPlugin_logic_onExecute_cmdSent <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        FpuSqrtPlugin_logic_onExecute_cmdSent <= 1'b0;
      end
      FpuSqrtPlugin_logic_onExecute_unscheduleRequest <= execute_lane0_ctrls_2_upIsCancel;
      if(execute_ctrl2_down_isReady) begin
        FpuSqrtPlugin_logic_onExecute_unscheduleRequest <= 1'b0;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_4) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      end
      decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= decode_ctrls_1_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l50_5) begin
        decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= 1'b0;
      end
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= execute_ctrl0_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_6) begin
        execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      execute_ctrl0_down_LANE_SEL_lane1_regNext <= execute_ctrl0_down_LANE_SEL_lane1;
      if(when_CtrlLaneApi_l50_7) begin
        execute_ctrl0_down_LANE_SEL_lane1_regNext <= 1'b0;
      end
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= execute_ctrl2_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_8) begin
        execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      execute_ctrl2_down_LANE_SEL_lane1_regNext <= execute_ctrl2_down_LANE_SEL_lane1;
      if(when_CtrlLaneApi_l50_9) begin
        execute_ctrl2_down_LANE_SEL_lane1_regNext <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))); // BtbPlugin.scala:L215
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L215
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[1]))); // BtbPlugin.scala:L215
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[1]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L215
            $finish;
          end
        `endif
      `endif
      if(fetch_logic_ctrls_1_up_isValid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l233) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      if(AlignerPlugin_logic_buffer_flushIt) begin
        AlignerPlugin_logic_buffer_mask <= 4'b0000;
        AlignerPlugin_logic_buffer_last <= 4'b0000;
      end
      if(DispatchPlugin_logic_slotsFeeds_doIt) begin
        DispatchPlugin_logic_slots_0_ctx_valid <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[0];
      end
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= TrapPlugin_logic_harts_0_interrupt_valid;
      PcPlugin_logic_harts_0_holdReg <= PcPlugin_logic_harts_0_holdComb;
      PcPlugin_logic_harts_0_self_state <= PcPlugin_logic_harts_0_output_payload_pc;
      PcPlugin_logic_harts_0_self_fault <= PcPlugin_logic_harts_0_output_payload_fault;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      if(PcPlugin_logic_harts_0_output_fire) begin
        PcPlugin_logic_harts_0_self_increment <= 1'b1;
        PcPlugin_logic_harts_0_self_state[2 : 1] <= 2'b00;
      end
      if(fetch_logic_ctrls_0_up_isFiring) begin
        PcPlugin_logic_harts_0_self_id <= (PcPlugin_logic_harts_0_self_id + 10'h001);
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))); // CsrAccessPlugin.scala:L136
        `else
          if(!(! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))) begin
            $display("FAILURE CsrAccessPlugin saw forbidden select && cancel request"); // CsrAccessPlugin.scala:L136
            $finish;
          end
        `endif
      `endif
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      if(CsrAccessPlugin_logic_flushPort_valid) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b1;
      end
      if(when_CsrAccessPlugin_l197) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      end
      CsrAccessPlugin_logic_fsm_inject_sampled <= execute_freeze_valid;
      if(when_CsrAccessPlugin_l346) begin
        PrefetcherRptPlugin_logic_csr_disable <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l346_1) begin
        PrivilegedPlugin_logic_harts_0_m_status_mpie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_status_mie <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= CsrAccessPlugin_bus_write_bits[17];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
      end
      if(when_CsrAccessPlugin_l346_2) begin
        PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= CsrAccessPlugin_bus_write_bits[31];
        PrivilegedPlugin_logic_harts_0_m_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l346_3) begin
        PrivilegedPlugin_logic_harts_0_m_ie_meie <= CsrAccessPlugin_bus_write_bits[11];
        PrivilegedPlugin_logic_harts_0_m_ie_mtie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_ie_msie <= CsrAccessPlugin_bus_write_bits[3];
      end
      if(when_CsrAccessPlugin_l346_4) begin
        FpuCsrPlugin_api_rm <= CsrAccessPlugin_bus_write_bits[7 : 5];
        FpuCsrPlugin_api_flags_NX <= _zz_FpuCsrPlugin_api_flags_NX[0];
        FpuCsrPlugin_api_flags_UF <= _zz_FpuCsrPlugin_api_flags_NX[1];
        FpuCsrPlugin_api_flags_OF <= _zz_FpuCsrPlugin_api_flags_NX[2];
        FpuCsrPlugin_api_flags_DZ <= _zz_FpuCsrPlugin_api_flags_NX[3];
        FpuCsrPlugin_api_flags_NV <= _zz_FpuCsrPlugin_api_flags_NX[4];
      end
      if(when_CsrAccessPlugin_l346_5) begin
        FpuCsrPlugin_api_rm <= CsrAccessPlugin_bus_write_bits[2 : 0];
      end
      if(when_CsrAccessPlugin_l346_6) begin
        FpuCsrPlugin_api_flags_NX <= _zz_FpuCsrPlugin_api_flags_NX_1[0];
        FpuCsrPlugin_api_flags_UF <= _zz_FpuCsrPlugin_api_flags_NX_1[1];
        FpuCsrPlugin_api_flags_OF <= _zz_FpuCsrPlugin_api_flags_NX_1[2];
        FpuCsrPlugin_api_flags_DZ <= _zz_FpuCsrPlugin_api_flags_NX_1[3];
        FpuCsrPlugin_api_flags_NV <= _zz_FpuCsrPlugin_api_flags_NX_1[4];
      end
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      CsrRamPlugin_logic_readLogic_ohReg <= (CsrRamPlugin_logic_readLogic_port_cmd_valid ? CsrRamPlugin_logic_readLogic_oh : 2'b00);
      CsrRamPlugin_logic_readLogic_busy <= CsrRamPlugin_logic_readLogic_port_cmd_valid;
      CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + _zz_CsrRamPlugin_logic_flush_counter);
      if(when_FpuFlagsWritebackPlugin_l96) begin
        if(FpuFlagsWritebackPlugin_logic_flagsOr_NV) begin
          FpuCsrPlugin_api_flags_NV <= 1'b1;
        end
        if(FpuFlagsWritebackPlugin_logic_flagsOr_DZ) begin
          FpuCsrPlugin_api_flags_DZ <= 1'b1;
        end
        if(FpuFlagsWritebackPlugin_logic_flagsOr_OF) begin
          FpuCsrPlugin_api_flags_OF <= 1'b1;
        end
        if(FpuFlagsWritebackPlugin_logic_flagsOr_UF) begin
          FpuCsrPlugin_api_flags_UF <= 1'b1;
        end
        if(FpuFlagsWritebackPlugin_logic_flagsOr_NX) begin
          FpuCsrPlugin_api_flags_NX <= 1'b1;
        end
      end
      if(when_RegFilePlugin_l132) begin
        integer_RegFilePlugin_logic_initalizer_counter <= (integer_RegFilePlugin_logic_initalizer_counter + 6'h01);
      end
      if(when_RegFilePlugin_l132_1) begin
        float_RegFilePlugin_logic_initalizer_counter <= (float_RegFilePlugin_logic_initalizer_counter + 6'h01);
      end
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
      if(fetch_logic_ctrls_1_up_forgetOne) begin
        fetch_logic_ctrls_1_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_0_down_isReady) begin
        fetch_logic_ctrls_1_up_valid <= fetch_logic_ctrls_0_down_isValid;
      end
      if(fetch_logic_ctrls_2_up_forgetOne) begin
        fetch_logic_ctrls_2_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_1_down_isReady) begin
        fetch_logic_ctrls_2_up_valid <= fetch_logic_ctrls_1_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_valid <= decode_ctrls_0_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_LANE_SEL_0 <= decode_ctrls_0_down_LANE_SEL_0;
        decode_ctrls_1_up_LANE_SEL_1 <= decode_ctrls_0_down_LANE_SEL_1;
      end
      if(when_DecodePipelinePlugin_l70) begin
        decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      end
      if(when_DecodePipelinePlugin_l70_1) begin
        decode_ctrls_1_up_LANE_SEL_1 <= 1'b0;
      end
      if(execute_ctrl0_down_isReady) begin
        execute_ctrl1_up_LANE_SEL_lane0 <= execute_ctrl0_down_LANE_SEL_lane0;
        execute_ctrl1_up_LANE_SEL_lane1 <= execute_ctrl0_down_LANE_SEL_lane1;
      end
      if(execute_ctrl1_down_isReady) begin
        execute_ctrl2_up_LANE_SEL_lane0 <= execute_ctrl1_down_LANE_SEL_lane0;
        execute_ctrl2_up_LANE_SEL_lane1 <= execute_ctrl1_down_LANE_SEL_lane1;
      end
      if(execute_ctrl2_down_isReady) begin
        execute_ctrl3_up_LANE_SEL_lane0 <= execute_ctrl2_down_LANE_SEL_lane0;
        execute_ctrl3_up_LANE_SEL_lane1 <= execute_ctrl2_down_LANE_SEL_lane1;
        execute_ctrl3_up_LsuL1_SEL_lane0 <= execute_ctrl2_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl3_down_isReady) begin
        execute_ctrl4_up_LANE_SEL_lane0 <= execute_ctrl3_down_LANE_SEL_lane0;
        execute_ctrl4_up_LANE_SEL_lane1 <= execute_ctrl3_down_LANE_SEL_lane1;
        execute_ctrl4_up_LsuL1_SEL_lane0 <= execute_ctrl3_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl4_down_isReady) begin
        execute_ctrl5_up_LANE_SEL_lane0 <= execute_ctrl4_down_LANE_SEL_lane0;
        execute_ctrl5_up_LANE_SEL_lane1 <= execute_ctrl4_down_LANE_SEL_lane1;
      end
      if(execute_ctrl5_down_isReady) begin
        execute_ctrl6_up_LANE_SEL_lane0 <= execute_ctrl5_down_LANE_SEL_lane0;
      end
      if(execute_ctrl6_down_isReady) begin
        execute_ctrl7_up_LANE_SEL_lane0 <= execute_ctrl6_down_LANE_SEL_lane0;
      end
      if(execute_ctrl7_down_isReady) begin
        execute_ctrl8_up_LANE_SEL_lane0 <= execute_ctrl7_down_LANE_SEL_lane0;
      end
      if(execute_ctrl8_down_isReady) begin
        execute_ctrl9_up_LANE_SEL_lane0 <= execute_ctrl8_down_LANE_SEL_lane0;
      end
      if(execute_ctrl9_down_isReady) begin
        execute_ctrl10_up_LANE_SEL_lane0 <= execute_ctrl9_down_LANE_SEL_lane0;
      end
      if(execute_ctrl10_down_isReady) begin
        execute_ctrl11_up_LANE_SEL_lane0 <= execute_ctrl10_down_LANE_SEL_lane0;
      end
      if(execute_ctrl11_down_isReady) begin
        execute_ctrl12_up_LANE_SEL_lane0 <= execute_ctrl11_down_LANE_SEL_lane0;
      end
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_stateNext;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_stateNext;
      case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
        TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
          TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
          if(!when_TrapPlugin_l409) begin
            case(TrapPlugin_logic_harts_0_trap_pending_state_code)
              4'b0000 : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert((! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)); // TrapPlugin.scala:L431
                  `else
                    if(!(! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)) begin
                      $display("FAILURE "); // TrapPlugin.scala:L431
                      $finish;
                    end
                  `endif
                `endif
              end
              4'b0001 : begin
              end
              4'b0010 : begin
              end
              4'b0100 : begin
              end
              4'b0101 : begin
              end
              4'b1000 : begin
              end
              4'b0110 : begin
              end
              default : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // TrapPlugin.scala:L482
                  `else
                    if(!1'b0) begin
                      $display("FAILURE Unexpected trap reason"); // TrapPlugin.scala:L482
                      $finish;
                    end
                  `endif
                `endif
              end
            endcase
          end
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
          case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= PrivilegedPlugin_logic_harts_0_m_status_mie;
              PrivilegedPlugin_logic_harts_0_m_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
          case(switch_TrapPlugin_l655)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mie <= PrivilegedPlugin_logic_harts_0_m_status_mpie;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        end
        default : begin
        end
      endcase
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_stateNext;
      case(CsrAccessPlugin_logic_fsm_stateReg)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
        end
        default : begin
          if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
            if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
              if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
                CsrAccessPlugin_logic_fsm_inject_unfreeze <= execute_freeze_valid;
              end
            end
          end
        end
      endcase
      case(CsrAccessPlugin_logic_fsm_stateNext)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
          CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b1;
        end
        default : begin
        end
      endcase
      BtbPlugin_logic_ras_ptr_pop <= BtbPlugin_logic_ras_ptr_pop_aheadValue;
    end
  end

  always @(posedge clk) begin
    LsuL1Plugin_logic_refill_slots_0_loadedCounter <= (LsuL1Plugin_logic_refill_slots_0_loadedCounter + ((LsuL1Plugin_logic_refill_slots_0_loaded && (! LsuL1Plugin_logic_refill_slots_0_loadedDone)) && (! execute_freeze_valid)));
    LsuL1Plugin_logic_refill_slots_1_loadedCounter <= (LsuL1Plugin_logic_refill_slots_1_loadedCounter + ((LsuL1Plugin_logic_refill_slots_1_loaded && (! LsuL1Plugin_logic_refill_slots_1_loadedDone)) && (! execute_freeze_valid)));
    if(LsuL1Plugin_logic_refill_slots_1_free) begin
      LsuL1Plugin_logic_refill_slots_0_priority[0] <= 1'b0;
    end
    if(when_LsuL1Plugin_l381) begin
      LsuL1Plugin_logic_refill_slots_0_address <= LsuL1Plugin_logic_refill_push_payload_address;
      LsuL1Plugin_logic_refill_slots_0_way <= LsuL1Plugin_logic_refill_push_payload_way;
      LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_priority <= 1'b1;
      LsuL1Plugin_logic_refill_slots_0_loadedCounter <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_victim <= LsuL1Plugin_logic_refill_push_payload_victim;
      LsuL1Plugin_logic_refill_slots_0_dirty <= LsuL1Plugin_logic_refill_push_payload_dirty;
    end
    if(LsuL1Plugin_logic_refill_slots_0_free) begin
      LsuL1Plugin_logic_refill_slots_1_priority[0] <= 1'b0;
    end
    if(when_LsuL1Plugin_l381_1) begin
      LsuL1Plugin_logic_refill_slots_1_address <= LsuL1Plugin_logic_refill_push_payload_address;
      LsuL1Plugin_logic_refill_slots_1_way <= LsuL1Plugin_logic_refill_push_payload_way;
      LsuL1Plugin_logic_refill_slots_1_cmdSent <= 1'b0;
      LsuL1Plugin_logic_refill_slots_1_priority <= 1'b1;
      LsuL1Plugin_logic_refill_slots_1_loadedCounter <= 1'b0;
      LsuL1Plugin_logic_refill_slots_1_victim <= LsuL1Plugin_logic_refill_push_payload_victim;
      LsuL1Plugin_logic_refill_slots_1_dirty <= LsuL1Plugin_logic_refill_push_payload_dirty;
    end
    if(LsuL1Plugin_logic_refill_read_arbiter_oh[0]) begin
      if(LsuL1Plugin_logic_bus_read_cmd_ready) begin
        LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      end
    end
    if(_zz_LsuL1Plugin_logic_refill_read_arbiter_sel) begin
      if(LsuL1Plugin_logic_bus_read_cmd_ready) begin
        LsuL1Plugin_logic_refill_slots_1_cmdSent <= 1'b1;
      end
    end
    LsuL1Plugin_logic_writeback_slots_0_timer_counter <= (LsuL1Plugin_logic_writeback_slots_0_timer_counter + ((! LsuL1Plugin_logic_writeback_slots_0_timer_done) && (! execute_freeze_valid)));
    LsuL1Plugin_logic_writeback_slots_1_timer_counter <= (LsuL1Plugin_logic_writeback_slots_1_timer_counter + ((! LsuL1Plugin_logic_writeback_slots_1_timer_done) && (! execute_freeze_valid)));
    if(LsuL1Plugin_logic_writeback_slots_1_free) begin
      LsuL1Plugin_logic_writeback_slots_0_priority[0] <= 1'b0;
    end
    if(when_LsuL1Plugin_l561) begin
      LsuL1Plugin_logic_writeback_slots_0_address <= LsuL1Plugin_logic_writeback_push_payload_address;
      LsuL1Plugin_logic_writeback_slots_0_way <= LsuL1Plugin_logic_writeback_push_payload_way;
      LsuL1Plugin_logic_writeback_slots_0_timer_counter <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_priority <= 1'b1;
      LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b0;
    end
    if(LsuL1Plugin_logic_writeback_slots_0_free) begin
      LsuL1Plugin_logic_writeback_slots_1_priority[0] <= 1'b0;
    end
    if(when_LsuL1Plugin_l561_1) begin
      LsuL1Plugin_logic_writeback_slots_1_address <= LsuL1Plugin_logic_writeback_push_payload_address;
      LsuL1Plugin_logic_writeback_slots_1_way <= LsuL1Plugin_logic_writeback_push_payload_way;
      LsuL1Plugin_logic_writeback_slots_1_timer_counter <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_writeCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_priority <= 1'b1;
      LsuL1Plugin_logic_writeback_slots_1_readCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_readRspDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_1_victimBufferReady <= 1'b0;
    end
    if(when_LsuL1Plugin_l605) begin
      if(LsuL1Plugin_logic_writeback_read_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b1;
      end
      if(_zz_LsuL1Plugin_logic_writeback_read_arbiter_sel) begin
        LsuL1Plugin_logic_writeback_slots_1_readCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_read_slotRead_valid) begin
      LsuL1Plugin_logic_refill_slots_0_victim[LsuL1Plugin_logic_writeback_read_slotRead_payload_id] <= 1'b0;
      LsuL1Plugin_logic_refill_slots_1_victim[LsuL1Plugin_logic_writeback_read_slotRead_payload_id] <= 1'b0;
    end
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_id <= LsuL1Plugin_logic_writeback_read_slotRead_payload_id;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last <= LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex <= LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way <= LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_id)
        1'b0 : begin
          LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b1;
        end
        default : begin
          LsuL1Plugin_logic_writeback_slots_1_victimBufferReady <= 1'b1;
        end
      endcase
      if(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last) begin
        case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_id)
          1'b0 : begin
            LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b1;
          end
          default : begin
            LsuL1Plugin_logic_writeback_slots_1_readRspDone <= 1'b1;
          end
        endcase
      end
    end
    if(when_LsuL1Plugin_l676) begin
      if(LsuL1Plugin_logic_writeback_write_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b1;
      end
      if(_zz_LsuL1Plugin_logic_writeback_write_arbiter_sel) begin
        LsuL1Plugin_logic_writeback_slots_1_writeCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_id <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_id;
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_address <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_last <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
    end
    if(PrefetcherRptPlugin_logic_pip2_node_0_isReady) begin
      PrefetcherRptPlugin_logic_pip2_node_1_CMD_address <= PrefetcherRptPlugin_logic_pip2_node_0_CMD_address;
      PrefetcherRptPlugin_logic_pip2_node_1_CMD_unique <= PrefetcherRptPlugin_logic_pip2_node_0_CMD_unique;
      PrefetcherRptPlugin_logic_pip2_node_1_CMD_from <= PrefetcherRptPlugin_logic_pip2_node_0_CMD_from;
      PrefetcherRptPlugin_logic_pip2_node_1_CMD_to <= PrefetcherRptPlugin_logic_pip2_node_0_CMD_to;
      PrefetcherRptPlugin_logic_pip2_node_1_CMD_stride <= PrefetcherRptPlugin_logic_pip2_node_0_CMD_stride;
      PrefetcherRptPlugin_logic_pip2_node_1_MUL <= PrefetcherRptPlugin_logic_pip2_node_0_MUL;
    end
    if(LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_ready) begin
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_last <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_last;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_write <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_write;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_id <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_id;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_address <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_address;
      LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_rData_fragment_data <= LsuL1Plugin_logic_bus_toWishbone_arbiter_serialized_payload_fragment_data;
    end
    if(when_FetchL1Plugin_l246) begin
      FetchL1Plugin_logic_refill_slots_0_priority[1] <= 1'b0;
    end
    if(when_FetchL1Plugin_l246_1) begin
      FetchL1Plugin_logic_refill_slots_1_priority[0] <= 1'b0;
    end
    if(when_FetchL1Plugin_l255) begin
      if(_zz_38) begin
        FetchL1Plugin_logic_refill_slots_0_address <= FetchL1Plugin_logic_refill_start_address;
        FetchL1Plugin_logic_refill_slots_0_isIo <= FetchL1Plugin_logic_refill_start_isIo;
        FetchL1Plugin_logic_refill_slots_0_wayToAllocate <= FetchL1Plugin_logic_refill_start_wayToAllocate;
        FetchL1Plugin_logic_refill_slots_0_priority <= {FetchL1Plugin_logic_refill_slots_1_valid,FetchL1Plugin_logic_refill_slots_0_valid};
      end
      if(_zz_when) begin
        FetchL1Plugin_logic_refill_slots_1_address <= FetchL1Plugin_logic_refill_start_address;
        FetchL1Plugin_logic_refill_slots_1_isIo <= FetchL1Plugin_logic_refill_start_isIo;
        FetchL1Plugin_logic_refill_slots_1_wayToAllocate <= FetchL1Plugin_logic_refill_start_wayToAllocate;
        FetchL1Plugin_logic_refill_slots_1_priority <= {FetchL1Plugin_logic_refill_slots_1_valid,FetchL1Plugin_logic_refill_slots_0_valid};
      end
    end
    if(when_FetchL1Plugin_l276) begin
      FetchL1Plugin_logic_refill_onCmd_lockedOh <= FetchL1Plugin_logic_refill_onCmd_propoedOh;
    end
    if(FetchL1Plugin_logic_bus_rsp_valid) begin
      FetchL1Plugin_logic_refill_onRsp_rspIdReg <= FetchL1Plugin_logic_bus_rsp_payload_id;
    end
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0 <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
    if(BtbPlugin_logic_ras_readIt) begin
      BtbPlugin_logic_ras_read <= BtbPlugin_logic_ras_mem_stack_spinal_port0;
    end
    FetchL1Plugin_logic_bus_cmd_payload_id_regNext <= FetchL1Plugin_logic_bus_cmd_payload_id;
    FetchL1WishbonePlugin_logic_bus_DAT_MISO_regNext <= FetchL1WishbonePlugin_logic_bus_DAT_MISO;
    FetchL1WishbonePlugin_logic_bus_ERR_regNext <= FetchL1WishbonePlugin_logic_bus_ERR;
    if(FpuAddSharedPlugin_logic_pip_node_0_isReady) begin
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mode;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_quiet <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_quiet;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_sign <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_sign;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_exponent;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mantissa <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs1_mantissa;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mode;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_quiet <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_quiet;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_sign <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_sign;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_exponent;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mantissa <= FpuAddSharedPlugin_logic_pip_node_0_inserter_rs2_mantissa;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FORMAT;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE <= FpuAddSharedPlugin_logic_pip_node_0_inserter_ROUNDMODE;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_RDN <= FpuAddSharedPlugin_logic_pip_node_0_inserter_RDN;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NX <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NX;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_UF <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_UF;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_OF <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_OF;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_DZ <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_DZ;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NV <= FpuAddSharedPlugin_logic_pip_node_0_inserter_FLAGS_NV;
      FpuAddSharedPlugin_logic_pip_node_1_Decode_UOP_ID <= FpuAddSharedPlugin_logic_pip_node_0_Decode_UOP_ID;
      FpuAddSharedPlugin_logic_pip_node_1_inserter_GROUP_OH <= FpuAddSharedPlugin_logic_pip_node_0_inserter_GROUP_OH;
      FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_absRs1Bigger <= FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_absRs1Bigger;
      FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_needSub <= FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_needSub;
      FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_passThrough <= FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_passThrough;
      FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_expDifAbsSat <= FpuAddSharedPlugin_logic_pip_node_0_adder_preShift_expDifAbsSat;
    end
    if(FpuAddSharedPlugin_logic_pip_node_1_isReady) begin
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mode;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_quiet <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_quiet;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_sign <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_sign;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_exponent;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mantissa <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs1_mantissa;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mode;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_quiet <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_quiet;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_sign <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_sign;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_exponent;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mantissa <= FpuAddSharedPlugin_logic_pip_node_1_inserter_rs2_mantissa;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FORMAT;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE <= FpuAddSharedPlugin_logic_pip_node_1_inserter_ROUNDMODE;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_RDN <= FpuAddSharedPlugin_logic_pip_node_1_inserter_RDN;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NX <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NX;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_UF <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_UF;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_OF <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_OF;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_DZ <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_DZ;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NV <= FpuAddSharedPlugin_logic_pip_node_1_inserter_FLAGS_NV;
      FpuAddSharedPlugin_logic_pip_node_2_Decode_UOP_ID <= FpuAddSharedPlugin_logic_pip_node_1_Decode_UOP_ID;
      FpuAddSharedPlugin_logic_pip_node_2_inserter_GROUP_OH <= FpuAddSharedPlugin_logic_pip_node_1_inserter_GROUP_OH;
      FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_needSub <= FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_needSub;
      FpuAddSharedPlugin_logic_pip_node_2_adder_preShift_passThrough <= FpuAddSharedPlugin_logic_pip_node_1_adder_preShift_passThrough;
      FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xySign <= FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xySign;
      FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xMantissa <= FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_xMantissa;
      FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_shifter <= FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_shifter;
      FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_yMantissa <= FpuAddSharedPlugin_logic_pip_node_1_adder_shifter_yMantissa;
      FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent <= _zz_FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xyExponent;
    end
    if(FpuAddSharedPlugin_logic_pip_node_2_isReady) begin
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mode;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_quiet <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_quiet;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_sign <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_sign;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_exponent;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mantissa <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs1_mantissa;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mode;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_quiet <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_quiet;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_sign <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_sign;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_exponent;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mantissa <= FpuAddSharedPlugin_logic_pip_node_2_inserter_rs2_mantissa;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FORMAT;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE <= FpuAddSharedPlugin_logic_pip_node_2_inserter_ROUNDMODE;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_RDN <= FpuAddSharedPlugin_logic_pip_node_2_inserter_RDN;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NX <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NX;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_UF <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_UF;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_OF <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_OF;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_DZ <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_DZ;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NV <= FpuAddSharedPlugin_logic_pip_node_2_inserter_FLAGS_NV;
      FpuAddSharedPlugin_logic_pip_node_3_Decode_UOP_ID <= FpuAddSharedPlugin_logic_pip_node_2_Decode_UOP_ID;
      FpuAddSharedPlugin_logic_pip_node_3_inserter_GROUP_OH <= FpuAddSharedPlugin_logic_pip_node_2_inserter_GROUP_OH;
      FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xySign <= FpuAddSharedPlugin_logic_pip_node_2_adder_shifter_xySign;
      FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent <= _zz_FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xyExponent;
      FpuAddSharedPlugin_logic_pip_node_3_adder_math_roundingScrap <= FpuAddSharedPlugin_logic_pip_node_2_adder_math_roundingScrap;
      FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa <= FpuAddSharedPlugin_logic_pip_node_2_adder_math_xyMantissa;
    end
    if(FpuAddSharedPlugin_logic_pip_node_3_isReady) begin
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mode <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mode;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_quiet <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_quiet;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_sign <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_sign;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_exponent;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs1_mantissa <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs1_mantissa;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mode <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mode;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_quiet <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_quiet;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_sign <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_sign;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_exponent <= _zz_FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_exponent;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_rs2_mantissa <= FpuAddSharedPlugin_logic_pip_node_3_inserter_rs2_mantissa;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FORMAT <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FORMAT;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_ROUNDMODE <= FpuAddSharedPlugin_logic_pip_node_3_inserter_ROUNDMODE;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_RDN <= FpuAddSharedPlugin_logic_pip_node_3_inserter_RDN;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NX <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NX;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_UF <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_UF;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_OF <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_OF;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_DZ <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_DZ;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_FLAGS_NV <= FpuAddSharedPlugin_logic_pip_node_3_inserter_FLAGS_NV;
      FpuAddSharedPlugin_logic_pip_node_4_Decode_UOP_ID <= FpuAddSharedPlugin_logic_pip_node_3_Decode_UOP_ID;
      FpuAddSharedPlugin_logic_pip_node_4_inserter_GROUP_OH <= FpuAddSharedPlugin_logic_pip_node_3_inserter_GROUP_OH;
      FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xySign <= FpuAddSharedPlugin_logic_pip_node_3_adder_shifter_xySign;
      FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent <= _zz_FpuAddSharedPlugin_logic_pip_node_4_adder_shifter_xyExponent;
      FpuAddSharedPlugin_logic_pip_node_4_adder_math_roundingScrap <= FpuAddSharedPlugin_logic_pip_node_3_adder_math_roundingScrap;
      FpuAddSharedPlugin_logic_pip_node_4_adder_math_xyMantissa <= FpuAddSharedPlugin_logic_pip_node_3_adder_math_xyMantissa;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_shift <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_shift;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceInfinity <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceInfinity;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceZero <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceZero;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_infinityNan <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_infinityNan;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_forceNan <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_forceNan;
      FpuAddSharedPlugin_logic_pip_node_4_adder_norm_xyMantissaZero <= FpuAddSharedPlugin_logic_pip_node_3_adder_norm_xyMantissaZero;
    end
    FpuUnpackerPlugin_logic_onUnpack_firstCycle <= 1'b0;
    if(when_FpuUnpackerPlugin_l165) begin
      FpuUnpackerPlugin_logic_onUnpack_firstCycle <= 1'b1;
    end
    early0_DivPlugin_logic_processing_divRevertResult <= ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ^ (execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 && (! execute_ctrl2_down_DivPlugin_REM_lane0))) && (! (((execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 == 32'h0) && execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0) && (! execute_ctrl2_down_DivPlugin_REM_lane0))));
    if(when_AlignerPlugin_l256) begin
      AlignerPlugin_logic_buffer_data <= fetch_logic_ctrls_2_down_Fetch_WORD;
      AlignerPlugin_logic_buffer_pc <= fetch_logic_ctrls_2_down_Fetch_WORD_PC;
      AlignerPlugin_logic_buffer_hm_Fetch_ID <= fetch_logic_ctrls_2_down_Fetch_ID;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3;
      AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
    end
    if(LsuPlugin_logic_storeBuffer_push_valid) begin
      if(_zz_when_3) begin
        LsuPlugin_logic_storeBuffer_slots_0_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_0_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_4) begin
        LsuPlugin_logic_storeBuffer_slots_1_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_1_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_5) begin
        LsuPlugin_logic_storeBuffer_slots_2_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_2_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_6) begin
        LsuPlugin_logic_storeBuffer_slots_3_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_3_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_7) begin
        LsuPlugin_logic_storeBuffer_slots_4_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_4_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_8) begin
        LsuPlugin_logic_storeBuffer_slots_5_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_5_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_9) begin
        LsuPlugin_logic_storeBuffer_slots_6_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_6_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
      if(_zz_when_10) begin
        LsuPlugin_logic_storeBuffer_slots_7_ptr <= LsuPlugin_logic_storeBuffer_ops_pushPtr;
        LsuPlugin_logic_storeBuffer_slots_7_tag <= LsuPlugin_logic_storeBuffer_push_payload_tag;
      end
    end
    if(LsuPlugin_logic_onAddress0_flush_port_fire) begin
      LsuPlugin_logic_flusher_cmdCounter <= (LsuPlugin_logic_flusher_cmdCounter + 7'h01);
    end
    if(LsuPlugin_logic_bus_rsp_toStream_ready) begin
      LsuPlugin_logic_bus_rsp_toStream_rData_error <= LsuPlugin_logic_bus_rsp_toStream_payload_error;
      LsuPlugin_logic_bus_rsp_toStream_rData_data <= LsuPlugin_logic_bus_rsp_toStream_payload_data;
    end
    LsuPlugin_logic_onCtrl_rva_srcBuffer <= execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0[31:0];
    LsuPlugin_logic_onCtrl_rva_aluBuffer <= LsuPlugin_logic_onCtrl_rva_alu_result;
    _zz_LsuPlugin_logic_onCtrl_rva_delay_0 <= (! execute_freeze_valid);
    _zz_LsuPlugin_logic_onCtrl_rva_delay_1 <= _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
    if(when_LsuPlugin_l698) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= (LsuPlugin_logic_onCtrl_rva_lrsc_age + 6'h01);
    end
    if(when_LsuPlugin_l705) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= 6'h0;
    end
    if(when_LsuPlugin_l709) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_address <= execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= 6'h0;
    end
    if(when_LsuPlugin_l905) begin
      LsuPlugin_logic_flusher_cmdCounter <= {1'd0, _zz_LsuPlugin_logic_flusher_cmdCounter};
    end
    if(when_LsuPlugin_l910) begin
      if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
        if(when_LsuPlugin_l913) begin
          if(when_LsuPlugin_l263) begin
            LsuPlugin_logic_storeBuffer_waitL1_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
          end
        end
      end
    end
    if(when_LsuPlugin_l949) begin
      if(when_LsuPlugin_l263_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    if(LsuPlugin_logic_storeBuffer_ops_pip_node_0_isReady) begin
      LsuPlugin_logic_storeBuffer_ops_pip_node_1_SB_PTR <= LsuPlugin_logic_storeBuffer_ops_pip_node_0_SB_PTR;
    end
    if(LsuPlugin_logic_storeBuffer_ops_pip_node_1_isReady) begin
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_SB_PTR <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_SB_PTR;
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_address <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_address;
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_data <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_data;
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_size <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_size;
      LsuPlugin_logic_storeBuffer_ops_pip_node_2_read_OPS_storeId <= LsuPlugin_logic_storeBuffer_ops_pip_node_1_read_OPS_storeId;
    end
    FpuPackerPlugin_logic_s1_subnormal_manShift <= _zz_FpuPackerPlugin_logic_s1_subnormal_manShift;
    FpuPackerPlugin_logic_s1_subnormal_manShifter <= _zz_FpuPackerPlugin_logic_s1_subnormal_manShifter_2[53 : 0];
    if(FpuPackerPlugin_logic_pip_node_0_isReady) begin
      FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode <= FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mode;
      FpuPackerPlugin_logic_pip_node_1_s0_VALUE_quiet <= FpuPackerPlugin_logic_pip_node_0_s0_VALUE_quiet;
      FpuPackerPlugin_logic_pip_node_1_s0_VALUE_sign <= FpuPackerPlugin_logic_pip_node_0_s0_VALUE_sign;
      FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent <= _zz_FpuPackerPlugin_logic_pip_node_1_s0_VALUE_exponent;
      FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mantissa <= FpuPackerPlugin_logic_pip_node_0_s0_VALUE_mantissa;
      FpuPackerPlugin_logic_pip_node_1_s0_FORMAT <= FpuPackerPlugin_logic_pip_node_0_s0_FORMAT;
      FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE <= FpuPackerPlugin_logic_pip_node_0_s0_ROUNDMODE;
      FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NX <= FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NX;
      FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_UF <= FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_UF;
      FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_OF <= FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_OF;
      FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_DZ <= FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_DZ;
      FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NV <= FpuPackerPlugin_logic_pip_node_0_s0_FLAGS_NV;
      FpuPackerPlugin_logic_pip_node_1_Decode_UOP_ID <= FpuPackerPlugin_logic_pip_node_0_Decode_UOP_ID;
      FpuPackerPlugin_logic_pip_node_1_s0_GROUP_OH <= FpuPackerPlugin_logic_pip_node_0_s0_GROUP_OH;
      FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL <= _zz_FpuPackerPlugin_logic_pip_node_1_s0_EXP_SUBNORMAL;
      FpuPackerPlugin_logic_pip_node_1_s0_subnormal_ENABLE <= FpuPackerPlugin_logic_pip_node_0_s0_subnormal_ENABLE;
    end
    if(FpuPackerPlugin_logic_pip_node_1_isReady) begin
      FpuPackerPlugin_logic_pip_node_2_s0_VALUE_mode <= FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mode;
      FpuPackerPlugin_logic_pip_node_2_s0_VALUE_quiet <= FpuPackerPlugin_logic_pip_node_1_s0_VALUE_quiet;
      FpuPackerPlugin_logic_pip_node_2_s0_VALUE_sign <= FpuPackerPlugin_logic_pip_node_1_s0_VALUE_sign;
      FpuPackerPlugin_logic_pip_node_2_s0_VALUE_exponent <= _zz_FpuPackerPlugin_logic_pip_node_2_s0_VALUE_exponent;
      FpuPackerPlugin_logic_s2_mr <= FpuPackerPlugin_logic_pip_node_1_s0_VALUE_mantissa;
      FpuPackerPlugin_logic_pip_node_2_s0_FORMAT <= FpuPackerPlugin_logic_pip_node_1_s0_FORMAT;
      FpuPackerPlugin_logic_pip_node_2_s0_ROUNDMODE <= FpuPackerPlugin_logic_pip_node_1_s0_ROUNDMODE;
      FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NX <= FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NX;
      FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_UF <= FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_UF;
      FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_OF <= FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_OF;
      FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_DZ <= FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_DZ;
      FpuPackerPlugin_logic_pip_node_2_s0_FLAGS_NV <= FpuPackerPlugin_logic_pip_node_1_s0_FLAGS_NV;
      FpuPackerPlugin_logic_pip_node_2_Decode_UOP_ID <= FpuPackerPlugin_logic_pip_node_1_Decode_UOP_ID;
      FpuPackerPlugin_logic_pip_node_2_s0_GROUP_OH <= FpuPackerPlugin_logic_pip_node_1_s0_GROUP_OH;
      FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL <= _zz_FpuPackerPlugin_logic_pip_node_2_s0_EXP_SUBNORMAL;
      FpuPackerPlugin_logic_pip_node_2_s0_subnormal_ENABLE <= FpuPackerPlugin_logic_pip_node_1_s0_subnormal_ENABLE;
      FpuPackerPlugin_logic_pip_node_2_s1_roundAdjusted <= FpuPackerPlugin_logic_pip_node_1_s1_roundAdjusted;
      FpuPackerPlugin_logic_pip_node_2_s1_manLsb <= FpuPackerPlugin_logic_pip_node_1_s1_manLsb;
      FpuPackerPlugin_logic_pip_node_2_s1_ROUNDING_INCR <= FpuPackerPlugin_logic_pip_node_1_s1_ROUNDING_INCR;
      FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT <= _zz_FpuPackerPlugin_logic_pip_node_2_s1_EXP_RESULT;
      FpuPackerPlugin_logic_pip_node_2_s1_MAN_RESULT <= FpuPackerPlugin_logic_pip_node_1_s1_MAN_RESULT;
    end
    if(LsuPlugin_logic_bus_cmd_ready) begin
      LsuPlugin_logic_bus_cmd_rData_write <= LsuPlugin_logic_bus_cmd_payload_write;
      LsuPlugin_logic_bus_cmd_rData_address <= LsuPlugin_logic_bus_cmd_payload_address;
      LsuPlugin_logic_bus_cmd_rData_data <= LsuPlugin_logic_bus_cmd_payload_data;
      LsuPlugin_logic_bus_cmd_rData_size <= LsuPlugin_logic_bus_cmd_payload_size;
      LsuPlugin_logic_bus_cmd_rData_mask <= LsuPlugin_logic_bus_cmd_payload_mask;
      LsuPlugin_logic_bus_cmd_rData_io <= LsuPlugin_logic_bus_cmd_payload_io;
      LsuPlugin_logic_bus_cmd_rData_fromHart <= LsuPlugin_logic_bus_cmd_payload_fromHart;
      LsuPlugin_logic_bus_cmd_rData_uopId <= LsuPlugin_logic_bus_cmd_payload_uopId;
    end
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_pc <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_pc;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_address <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_address;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_load <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_load;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_store <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_store;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_trap <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_trap;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_io <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_io;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_prefetchFailed <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_prefetchFailed;
    PrefetcherRptPlugin_logic_pip_node_1_PROBE_miss <= PrefetcherRptPlugin_logic_pip_node_0_PROBE_miss;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_valid <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_valid;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_address <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_address;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_tag <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_tag;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_address <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_address;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_stride <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_stride;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_score <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_score;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_advance <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_advance;
    PrefetcherRptPlugin_logic_pip_node_1_onRead0_WRITTEN_payload_data_missed <= PrefetcherRptPlugin_logic_pip_node_0_onRead0_WRITTEN_payload_data_missed;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_pc <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_pc;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_address <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_address;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_load <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_load;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_store <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_store;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_trap <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_trap;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_io <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_io;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_prefetchFailed <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_prefetchFailed;
    PrefetcherRptPlugin_logic_pip_node_2_PROBE_miss <= PrefetcherRptPlugin_logic_pip_node_1_PROBE_miss;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_tag <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_tag;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_address <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_address;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_stride <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_stride;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_score <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_score;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_advance <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_advance;
    PrefetcherRptPlugin_logic_pip_node_2_ENTRY_missed <= PrefetcherRptPlugin_logic_pip_node_1_ENTRY_missed;
    PrefetcherRptPlugin_logic_pip_node_2_TAG_HIT <= PrefetcherRptPlugin_logic_pip_node_1_TAG_HIT;
    PrefetcherRptPlugin_logic_pip_node_2_STRIDE_EXTENDED <= PrefetcherRptPlugin_logic_pip_node_1_STRIDE_EXTENDED;
    PrefetcherRptPlugin_logic_pip_node_2_NEW_BLOCK <= PrefetcherRptPlugin_logic_pip_node_1_NEW_BLOCK;
    if(late0_BranchPlugin_logic_jumpLogic_learn_ready) begin
      late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice <= late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget <= late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_taken <= late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong <= late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget <= late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_history <= late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId <= late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
    end
    if(late1_BranchPlugin_logic_jumpLogic_learn_ready) begin
      late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice <= late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget <= late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_taken <= late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong <= late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget <= late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_history <= late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId <= late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
    end
    if(when_FpuUnpackerPlugin_l251) begin
      FpuUnpack_RS1_normalizer_exponent <= _zz_FpuUnpack_RS1_normalizer_exponent;
      FpuUnpack_RS1_normalizer_mantissa <= FpuUnpackerPlugin_logic_unpacker_results_0_payload_data;
    end
    if(when_FpuUnpackerPlugin_l251_1) begin
      FpuUnpack_RS2_normalizer_exponent <= _zz_FpuUnpack_RS2_normalizer_exponent;
      FpuUnpack_RS2_normalizer_mantissa <= FpuUnpackerPlugin_logic_unpacker_results_0_payload_data;
    end
    if(when_FpuUnpackerPlugin_l251_2) begin
      FpuUnpack_RS3_normalizer_exponent <= _zz_FpuUnpack_RS3_normalizer_exponent;
      FpuUnpack_RS3_normalizer_mantissa <= FpuUnpackerPlugin_logic_unpacker_results_0_payload_data;
    end
    if(FpuUnpackerPlugin_logic_unpacker_results_1_valid) begin
      FpuUnpackerPlugin_logic_onCvt_fsmResult_shift <= FpuUnpackerPlugin_logic_unpacker_results_1_payload_shift;
      FpuUnpackerPlugin_logic_onCvt_fsmResult_data <= FpuUnpackerPlugin_logic_unpacker_results_1_payload_data;
    end
    FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data <= FpuUnpackerPlugin_logic_unpacker_node_0_input_args_data;
    FpuUnpackerPlugin_logic_unpacker_node_1_input_source <= FpuUnpackerPlugin_logic_unpacker_node_0_input_source;
    FpuUnpackerPlugin_logic_unpacker_node_2_input_args_data <= FpuUnpackerPlugin_logic_unpacker_node_1_input_args_data;
    FpuUnpackerPlugin_logic_unpacker_node_2_input_source <= FpuUnpackerPlugin_logic_unpacker_node_1_input_source;
    FpuUnpackerPlugin_logic_unpacker_node_2_setup_shiftBy <= FpuUnpackerPlugin_logic_unpacker_node_1_setup_shiftBy;
    FpuF2iPlugin_logic_onResult_inverter <= ((execute_ctrl4_down_FpuF2iPlugin_logic_onShift_resign_lane0 ? (~ FpuF2iPlugin_logic_onResult_unsigned) : FpuF2iPlugin_logic_onResult_unsigned) + _zz_FpuF2iPlugin_logic_onResult_inverter);
    _zz_FpuDivPlugin_logic_onExecute_exponent <= _zz__zz_FpuDivPlugin_logic_onExecute_exponent;
    if(DispatchPlugin_logic_slotsFeeds_doIt) begin
      DispatchPlugin_logic_slots_0_ctx_laneLayerHits <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[4 : 1];
      DispatchPlugin_logic_slots_0_ctx_uop <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[36 : 5];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[0];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[32 : 1];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[36 : 33];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[40 : 37];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[1 : 0];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[3 : 2];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[5 : 4];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[7 : 6];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[60 : 49];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[61];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[62];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[63];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[64];
      DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[65 : 65];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_2 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[66];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_6 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[67];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_5 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[68];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[69];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_9 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[70];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_2 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[71];
      DispatchPlugin_logic_slots_0_ctx_hm_FpuPackerPlugin_RESERVED_ON_early0_AT_3 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[72];
      DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[73];
      DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[74];
      DispatchPlugin_logic_slots_0_ctx_hm_PC <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[106 : 75];
      DispatchPlugin_logic_slots_0_ctx_hm_TRAP <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[107];
      DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[123 : 108];
      DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[124];
      DispatchPlugin_logic_slots_0_ctx_hm_RS1_RFID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[125 : 125];
      DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[130 : 126];
      DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[131];
      DispatchPlugin_logic_slots_0_ctx_hm_RS2_RFID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[132 : 132];
      DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[137 : 133];
      DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[138];
      DispatchPlugin_logic_slots_0_ctx_hm_RD_RFID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[139 : 139];
      DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[144 : 140];
      DispatchPlugin_logic_slots_0_ctx_hm_RS3_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[145];
      DispatchPlugin_logic_slots_0_ctx_hm_RS3_RFID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[146 : 146];
      DispatchPlugin_logic_slots_0_ctx_hm_RS3_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[151 : 147];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[152];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[153];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[154];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[155];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_2_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[156];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[157];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[158];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[159];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[160];
    end
    if(TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_state_exception <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
      TrapPlugin_logic_harts_0_trap_pending_state_tval <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
      TrapPlugin_logic_harts_0_trap_pending_state_code <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
      TrapPlugin_logic_harts_0_trap_pending_state_arg <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
    end
    if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_pc <= ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? execute_ctrl4_down_PC_lane0 : 32'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? execute_ctrl4_down_PC_lane1 : 32'h0));
      TrapPlugin_logic_harts_0_trap_pending_history <= ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 : 12'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1 : 12'h0));
      TrapPlugin_logic_harts_0_trap_pending_slices <= (_zz_TrapPlugin_logic_harts_0_trap_pending_slices + 2'b01);
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid <= TrapPlugin_logic_harts_0_interrupt_valid;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code <= TrapPlugin_logic_harts_0_interrupt_code;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege <= TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
    end
    TrapPlugin_logic_harts_0_trap_fsm_jumpTarget <= (TrapPlugin_logic_harts_0_trap_pending_pc + _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget);
    if(when_TrapPlugin_l556) begin
      TrapPlugin_logic_harts_0_trap_fsm_readed <= TrapPlugin_logic_harts_0_crsPorts_read_data;
    end
    CsrAccessPlugin_logic_fsm_interface_read <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrRead);
    CsrAccessPlugin_logic_fsm_interface_write <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrWrite);
    CsrAccessPlugin_logic_fsm_inject_trapReg <= CsrAccessPlugin_logic_fsm_inject_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapReg <= CsrAccessPlugin_bus_decode_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg <= CsrAccessPlugin_bus_decode_trapCode;
    CsrAccessPlugin_logic_fsm_interface_onWriteBits <= CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(fetch_logic_ctrls_0_down_isReady) begin
      fetch_logic_ctrls_1_up_Fetch_WORD_PC <= fetch_logic_ctrls_0_down_Fetch_WORD_PC;
      fetch_logic_ctrls_1_up_Fetch_PC_FAULT <= fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_1_up_Fetch_ID <= fetch_logic_ctrls_0_down_Fetch_ID;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH <= fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
      fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3;
      fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS <= fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
    end
    if(fetch_logic_ctrls_1_down_isReady) begin
      fetch_logic_ctrls_2_up_Fetch_WORD_PC <= fetch_logic_ctrls_1_down_Fetch_WORD_PC;
      fetch_logic_ctrls_2_up_Fetch_PC_FAULT <= fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_2_up_Fetch_ID <= fetch_logic_ctrls_1_down_Fetch_ID;
      fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
      fetch_logic_ctrls_2_up_MMU_TRANSLATED <= fetch_logic_ctrls_1_down_MMU_TRANSLATED;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_SLICE <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_SLICE;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
      fetch_logic_ctrls_2_up_MMU_REFILL <= fetch_logic_ctrls_1_down_MMU_REFILL;
      fetch_logic_ctrls_2_up_MMU_HAZARD <= fetch_logic_ctrls_1_down_MMU_HAZARD;
      fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE <= fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
      fetch_logic_ctrls_2_up_MMU_PAGE_FAULT <= fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
      fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT <= fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
      fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION <= fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
    end
    if(decode_ctrls_0_down_isReady) begin
      decode_ctrls_1_up_Decode_INSTRUCTION_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_0;
      decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0 <= decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
      decode_ctrls_1_up_PC_0 <= decode_ctrls_0_down_PC_0;
      decode_ctrls_1_up_Decode_DOP_ID_0 <= decode_ctrls_0_down_Decode_DOP_ID_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3;
      decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0 <= decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
      decode_ctrls_1_up_TRAP_0 <= decode_ctrls_0_down_TRAP_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
      decode_ctrls_1_up_Prediction_ALIGN_REDO_0 <= decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_1 <= decode_ctrls_0_down_Decode_INSTRUCTION_1;
      decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1 <= decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1;
      decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1 <= decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1;
      decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1 <= decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1;
      decode_ctrls_1_up_PC_1 <= decode_ctrls_0_down_PC_1;
      decode_ctrls_1_up_Decode_DOP_ID_1 <= decode_ctrls_0_down_Decode_DOP_ID_1;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3;
      decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1 <= decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1;
      decode_ctrls_1_up_TRAP_1 <= decode_ctrls_0_down_TRAP_1;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1;
      decode_ctrls_1_up_Prediction_ALIGN_REDO_1 <= decode_ctrls_0_down_Prediction_ALIGN_REDO_1;
    end
    if(execute_ctrl0_down_isReady) begin
      execute_ctrl1_up_Decode_UOP_lane0 <= execute_ctrl0_down_Decode_UOP_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 <= execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
      execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl1_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl0_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl1_up_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0 <= execute_ctrl0_down_FpuPackerPlugin_RESERVED_ON_early0_AT_3_lane0;
      execute_ctrl1_up_PC_lane0 <= execute_ctrl0_down_PC_lane0;
      execute_ctrl1_up_TRAP_lane0 <= execute_ctrl0_down_TRAP_lane0;
      execute_ctrl1_up_Decode_UOP_ID_lane0 <= execute_ctrl0_down_Decode_UOP_ID_lane0;
      execute_ctrl1_up_RS1_ENABLE_lane0 <= execute_ctrl0_down_RS1_ENABLE_lane0;
      execute_ctrl1_up_RS1_RFID_lane0 <= execute_ctrl0_down_RS1_RFID_lane0;
      execute_ctrl1_up_RS1_PHYS_lane0 <= execute_ctrl0_down_RS1_PHYS_lane0;
      execute_ctrl1_up_RS2_ENABLE_lane0 <= execute_ctrl0_down_RS2_ENABLE_lane0;
      execute_ctrl1_up_RS2_RFID_lane0 <= execute_ctrl0_down_RS2_RFID_lane0;
      execute_ctrl1_up_RS2_PHYS_lane0 <= execute_ctrl0_down_RS2_PHYS_lane0;
      execute_ctrl1_up_RD_ENABLE_lane0 <= execute_ctrl0_down_RD_ENABLE_lane0;
      execute_ctrl1_up_RD_RFID_lane0 <= execute_ctrl0_down_RD_RFID_lane0;
      execute_ctrl1_up_RD_PHYS_lane0 <= execute_ctrl0_down_RD_PHYS_lane0;
      execute_ctrl1_up_RS3_ENABLE_lane0 <= execute_ctrl0_down_RS3_ENABLE_lane0;
      execute_ctrl1_up_RS3_RFID_lane0 <= execute_ctrl0_down_RS3_RFID_lane0;
      execute_ctrl1_up_RS3_PHYS_lane0 <= execute_ctrl0_down_RS3_PHYS_lane0;
      execute_ctrl1_up_LANE_AGE_lane0 <= execute_ctrl0_down_LANE_AGE_lane0;
      execute_ctrl1_up_COMPLETED_lane0 <= execute_ctrl0_down_COMPLETED_lane0;
      execute_ctrl1_up_lane0_LAYER_SEL_lane0 <= execute_ctrl0_down_lane0_LAYER_SEL_lane0;
      execute_ctrl1_up_Decode_UOP_lane1 <= execute_ctrl0_down_Decode_UOP_lane1;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1 <= execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1;
      execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      execute_ctrl1_up_PC_lane1 <= execute_ctrl0_down_PC_lane1;
      execute_ctrl1_up_TRAP_lane1 <= execute_ctrl0_down_TRAP_lane1;
      execute_ctrl1_up_Decode_UOP_ID_lane1 <= execute_ctrl0_down_Decode_UOP_ID_lane1;
      execute_ctrl1_up_RS1_RFID_lane1 <= execute_ctrl0_down_RS1_RFID_lane1;
      execute_ctrl1_up_RS1_PHYS_lane1 <= execute_ctrl0_down_RS1_PHYS_lane1;
      execute_ctrl1_up_RS2_RFID_lane1 <= execute_ctrl0_down_RS2_RFID_lane1;
      execute_ctrl1_up_RS2_PHYS_lane1 <= execute_ctrl0_down_RS2_PHYS_lane1;
      execute_ctrl1_up_RD_ENABLE_lane1 <= execute_ctrl0_down_RD_ENABLE_lane1;
      execute_ctrl1_up_RD_RFID_lane1 <= execute_ctrl0_down_RD_RFID_lane1;
      execute_ctrl1_up_RD_PHYS_lane1 <= execute_ctrl0_down_RD_PHYS_lane1;
      execute_ctrl1_up_LANE_AGE_lane1 <= execute_ctrl0_down_LANE_AGE_lane1;
      execute_ctrl1_up_COMPLETED_lane1 <= execute_ctrl0_down_COMPLETED_lane1;
      execute_ctrl1_up_lane1_LAYER_SEL_lane1 <= execute_ctrl0_down_lane1_LAYER_SEL_lane1;
      execute_ctrl1_up_AguPlugin_SIZE_lane0 <= execute_ctrl0_down_AguPlugin_SIZE_lane0;
    end
    if(execute_ctrl1_down_isReady) begin
      execute_ctrl2_up_Decode_UOP_lane0 <= execute_ctrl1_down_Decode_UOP_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 <= execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
      execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl2_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl1_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl2_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl1_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl2_up_PC_lane0 <= execute_ctrl1_down_PC_lane0;
      execute_ctrl2_up_TRAP_lane0 <= execute_ctrl1_down_TRAP_lane0;
      execute_ctrl2_up_Decode_UOP_ID_lane0 <= execute_ctrl1_down_Decode_UOP_ID_lane0;
      execute_ctrl2_up_RS1_ENABLE_lane0 <= execute_ctrl1_down_RS1_ENABLE_lane0;
      execute_ctrl2_up_RS1_RFID_lane0 <= execute_ctrl1_down_RS1_RFID_lane0;
      execute_ctrl2_up_RS1_PHYS_lane0 <= execute_ctrl1_down_RS1_PHYS_lane0;
      execute_ctrl2_up_RS2_ENABLE_lane0 <= execute_ctrl1_down_RS2_ENABLE_lane0;
      execute_ctrl2_up_RS2_RFID_lane0 <= execute_ctrl1_down_RS2_RFID_lane0;
      execute_ctrl2_up_RS2_PHYS_lane0 <= execute_ctrl1_down_RS2_PHYS_lane0;
      execute_ctrl2_up_RD_ENABLE_lane0 <= execute_ctrl1_down_RD_ENABLE_lane0;
      execute_ctrl2_up_RD_RFID_lane0 <= execute_ctrl1_down_RD_RFID_lane0;
      execute_ctrl2_up_RD_PHYS_lane0 <= execute_ctrl1_down_RD_PHYS_lane0;
      execute_ctrl2_up_RS3_ENABLE_lane0 <= execute_ctrl1_down_RS3_ENABLE_lane0;
      execute_ctrl2_up_RS3_RFID_lane0 <= execute_ctrl1_down_RS3_RFID_lane0;
      execute_ctrl2_up_LANE_AGE_lane0 <= execute_ctrl1_down_LANE_AGE_lane0;
      execute_ctrl2_up_COMPLETED_lane0 <= execute_ctrl1_down_COMPLETED_lane0;
      execute_ctrl2_up_Decode_UOP_lane1 <= execute_ctrl1_down_Decode_UOP_lane1;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1 <= execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1;
      execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      execute_ctrl2_up_PC_lane1 <= execute_ctrl1_down_PC_lane1;
      execute_ctrl2_up_TRAP_lane1 <= execute_ctrl1_down_TRAP_lane1;
      execute_ctrl2_up_Decode_UOP_ID_lane1 <= execute_ctrl1_down_Decode_UOP_ID_lane1;
      execute_ctrl2_up_RS1_RFID_lane1 <= execute_ctrl1_down_RS1_RFID_lane1;
      execute_ctrl2_up_RS1_PHYS_lane1 <= execute_ctrl1_down_RS1_PHYS_lane1;
      execute_ctrl2_up_RS2_RFID_lane1 <= execute_ctrl1_down_RS2_RFID_lane1;
      execute_ctrl2_up_RS2_PHYS_lane1 <= execute_ctrl1_down_RS2_PHYS_lane1;
      execute_ctrl2_up_RD_ENABLE_lane1 <= execute_ctrl1_down_RD_ENABLE_lane1;
      execute_ctrl2_up_RD_RFID_lane1 <= execute_ctrl1_down_RD_RFID_lane1;
      execute_ctrl2_up_RD_PHYS_lane1 <= execute_ctrl1_down_RD_PHYS_lane1;
      execute_ctrl2_up_LANE_AGE_lane1 <= execute_ctrl1_down_LANE_AGE_lane1;
      execute_ctrl2_up_COMPLETED_lane1 <= execute_ctrl1_down_COMPLETED_lane1;
      execute_ctrl2_up_AguPlugin_SIZE_lane0 <= execute_ctrl1_down_AguPlugin_SIZE_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
      execute_ctrl2_up_integer_RS1_lane0 <= execute_ctrl1_down_integer_RS1_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
      execute_ctrl2_up_integer_RS2_lane0 <= execute_ctrl1_down_integer_RS2_lane0;
      execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1 <= execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
      execute_ctrl2_up_integer_RS1_lane1 <= execute_ctrl1_down_integer_RS1_lane1;
      execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1 <= execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
      execute_ctrl2_up_integer_RS2_lane1 <= execute_ctrl1_down_integer_RS2_lane1;
      execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0 <= execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
      execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1 <= execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
      execute_ctrl2_up_float_RS1_lane0 <= execute_ctrl1_down_float_RS1_lane0;
      execute_ctrl2_up_float_RS2_lane0 <= execute_ctrl1_down_float_RS2_lane0;
      execute_ctrl2_up_float_RS3_lane0 <= execute_ctrl1_down_float_RS3_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl2_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl2_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl2_up_early0_EnvPlugin_SEL_lane0 <= execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
      execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0 <= execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
      execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl2_up_late0_BranchPlugin_SEL_lane0 <= execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
      execute_ctrl2_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl2_up_FpuCsrPlugin_DIRTY_lane0 <= execute_ctrl1_down_FpuCsrPlugin_DIRTY_lane0;
      execute_ctrl2_up_FpuClassPlugin_SEL_lane0 <= execute_ctrl1_down_FpuClassPlugin_SEL_lane0;
      execute_ctrl2_up_FpuCmpPlugin_SEL_FLOAT_lane0 <= execute_ctrl1_down_FpuCmpPlugin_SEL_FLOAT_lane0;
      execute_ctrl2_up_FpuCmpPlugin_SEL_CMP_lane0 <= execute_ctrl1_down_FpuCmpPlugin_SEL_CMP_lane0;
      execute_ctrl2_up_FpuF2iPlugin_SEL_lane0 <= execute_ctrl1_down_FpuF2iPlugin_SEL_lane0;
      execute_ctrl2_up_FpuMvPlugin_SEL_FLOAT_lane0 <= execute_ctrl1_down_FpuMvPlugin_SEL_FLOAT_lane0;
      execute_ctrl2_up_FpuMvPlugin_SEL_INT_lane0 <= execute_ctrl1_down_FpuMvPlugin_SEL_INT_lane0;
      execute_ctrl2_up_AguPlugin_SEL_lane0 <= execute_ctrl1_down_AguPlugin_SEL_lane0;
      execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl2_up_FpuAddPlugin_SEL_lane0 <= execute_ctrl1_down_FpuAddPlugin_SEL_lane0;
      execute_ctrl2_up_FpuMulPlugin_SEL_lane0 <= execute_ctrl1_down_FpuMulPlugin_SEL_lane0;
      execute_ctrl2_up_FpuSqrtPlugin_SEL_lane0 <= execute_ctrl1_down_FpuSqrtPlugin_SEL_lane0;
      execute_ctrl2_up_FpuXxPlugin_SEL_lane0 <= execute_ctrl1_down_FpuXxPlugin_SEL_lane0;
      execute_ctrl2_up_FpuDivPlugin_SEL_lane0 <= execute_ctrl1_down_FpuDivPlugin_SEL_lane0;
      execute_ctrl2_up_FpuUnpackerPlugin_SEL_I2F_lane0 <= execute_ctrl1_down_FpuUnpackerPlugin_SEL_I2F_lane0;
      execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl2_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl1_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl2_up_COMPLETION_AT_4_lane0 <= execute_ctrl1_down_COMPLETION_AT_4_lane0;
      execute_ctrl2_up_COMPLETION_AT_7_lane0 <= execute_ctrl1_down_COMPLETION_AT_7_lane0;
      execute_ctrl2_up_COMPLETION_AT_11_lane0 <= execute_ctrl1_down_COMPLETION_AT_11_lane0;
      execute_ctrl2_up_COMPLETION_AT_3_lane0 <= execute_ctrl1_down_COMPLETION_AT_3_lane0;
      execute_ctrl2_up_COMPLETION_AT_5_lane0 <= execute_ctrl1_down_COMPLETION_AT_5_lane0;
      execute_ctrl2_up_COMPLETION_AT_8_lane0 <= execute_ctrl1_down_COMPLETION_AT_8_lane0;
      execute_ctrl2_up_COMPLETION_AT_2_lane0 <= execute_ctrl1_down_COMPLETION_AT_2_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_6_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_6_ENABLE_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl2_up_SrcStageables_REVERT_lane0 <= execute_ctrl1_down_SrcStageables_REVERT_lane0;
      execute_ctrl2_up_SrcStageables_ZERO_lane0 <= execute_ctrl1_down_SrcStageables_ZERO_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl2_up_BYPASSED_AT_3_lane0 <= execute_ctrl1_down_BYPASSED_AT_3_lane0;
      execute_ctrl2_up_BYPASSED_AT_4_lane0 <= execute_ctrl1_down_BYPASSED_AT_4_lane0;
      execute_ctrl2_up_BYPASSED_AT_5_lane0 <= execute_ctrl1_down_BYPASSED_AT_5_lane0;
      execute_ctrl2_up_BYPASSED_AT_6_lane0 <= execute_ctrl1_down_BYPASSED_AT_6_lane0;
      execute_ctrl2_up_BYPASSED_AT_7_lane0 <= execute_ctrl1_down_BYPASSED_AT_7_lane0;
      execute_ctrl2_up_BYPASSED_AT_8_lane0 <= execute_ctrl1_down_BYPASSED_AT_8_lane0;
      execute_ctrl2_up_BYPASSED_AT_9_lane0 <= execute_ctrl1_down_BYPASSED_AT_9_lane0;
      execute_ctrl2_up_BYPASSED_AT_10_lane0 <= execute_ctrl1_down_BYPASSED_AT_10_lane0;
      execute_ctrl2_up_SrcStageables_UNSIGNED_lane0 <= execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
      execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl2_up_MulPlugin_HIGH_lane0 <= execute_ctrl1_down_MulPlugin_HIGH_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
      execute_ctrl2_up_DivPlugin_REM_lane0 <= execute_ctrl1_down_DivPlugin_REM_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
      execute_ctrl2_up_FpuUtils_FORMAT_lane0 <= execute_ctrl1_down_FpuUtils_FORMAT_lane0;
      execute_ctrl2_up_FpuCmpPlugin_FLOAT_OP_lane0 <= execute_ctrl1_down_FpuCmpPlugin_FLOAT_OP_lane0;
      execute_ctrl2_up_FpuCmpPlugin_INVERT_lane0 <= execute_ctrl1_down_FpuCmpPlugin_INVERT_lane0;
      execute_ctrl2_up_FpuCmpPlugin_SGNJ_RS1_lane0 <= execute_ctrl1_down_FpuCmpPlugin_SGNJ_RS1_lane0;
      execute_ctrl2_up_FpuCmpPlugin_LESS_lane0 <= execute_ctrl1_down_FpuCmpPlugin_LESS_lane0;
      execute_ctrl2_up_FpuCmpPlugin_EQUAL_lane0 <= execute_ctrl1_down_FpuCmpPlugin_EQUAL_lane0;
      execute_ctrl2_up_AguPlugin_LOAD_lane0 <= execute_ctrl1_down_AguPlugin_LOAD_lane0;
      execute_ctrl2_up_AguPlugin_STORE_lane0 <= execute_ctrl1_down_AguPlugin_STORE_lane0;
      execute_ctrl2_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl2_up_AguPlugin_FLOAT_lane0 <= execute_ctrl1_down_AguPlugin_FLOAT_lane0;
      execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl2_up_early0_EnvPlugin_OP_lane0 <= execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
      execute_ctrl2_up_FpuAddPlugin_SUB_lane0 <= execute_ctrl1_down_FpuAddPlugin_SUB_lane0;
      execute_ctrl2_up_FpuMulPlugin_FMA_lane0 <= execute_ctrl1_down_FpuMulPlugin_FMA_lane0;
      execute_ctrl2_up_FpuMulPlugin_SUB1_lane0 <= execute_ctrl1_down_FpuMulPlugin_SUB1_lane0;
      execute_ctrl2_up_FpuMulPlugin_SUB2_lane0 <= execute_ctrl1_down_FpuMulPlugin_SUB2_lane0;
      execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0 <= execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
      execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0 <= execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
      execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1 <= execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
      execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1 <= execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
      execute_ctrl2_up_early1_BranchPlugin_SEL_lane1 <= execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
      execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1 <= execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
      execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1 <= execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
      execute_ctrl2_up_late1_BranchPlugin_SEL_lane1 <= execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
      execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      execute_ctrl2_up_COMPLETION_AT_2_lane1 <= execute_ctrl1_down_COMPLETION_AT_2_lane1;
      execute_ctrl2_up_COMPLETION_AT_4_lane1 <= execute_ctrl1_down_COMPLETION_AT_4_lane1;
      execute_ctrl2_up_lane1_logic_completions_onCtrl_0_ENABLE_lane1 <= execute_ctrl1_down_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
      execute_ctrl2_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1 <= execute_ctrl1_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
      execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1 <= execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
      execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1 <= execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
      execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      execute_ctrl2_up_SrcStageables_REVERT_lane1 <= execute_ctrl1_down_SrcStageables_REVERT_lane1;
      execute_ctrl2_up_SrcStageables_ZERO_lane1 <= execute_ctrl1_down_SrcStageables_ZERO_lane1;
      execute_ctrl2_up_BYPASSED_AT_3_lane1 <= execute_ctrl1_down_BYPASSED_AT_3_lane1;
      execute_ctrl2_up_SrcStageables_UNSIGNED_lane1 <= execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
      execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1 <= execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
      execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1 <= execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
      execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1 <= execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
      execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1 <= execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
      execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1 <= execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
    end
    if(execute_ctrl2_down_isReady) begin
      execute_ctrl3_up_Decode_UOP_lane0 <= execute_ctrl2_down_Decode_UOP_lane0;
      execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 <= execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
      execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl3_up_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0 <= execute_ctrl2_down_FpuAddSharedPlugin_RESERVED_ON_early0_AT_5_lane0;
      execute_ctrl3_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl2_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl3_up_PC_lane0 <= execute_ctrl2_down_PC_lane0;
      execute_ctrl3_up_TRAP_lane0 <= execute_ctrl2_down_TRAP_lane0;
      execute_ctrl3_up_Decode_UOP_ID_lane0 <= execute_ctrl2_down_Decode_UOP_ID_lane0;
      execute_ctrl3_up_RS1_RFID_lane0 <= execute_ctrl2_down_RS1_RFID_lane0;
      execute_ctrl3_up_RS1_PHYS_lane0 <= execute_ctrl2_down_RS1_PHYS_lane0;
      execute_ctrl3_up_RS2_RFID_lane0 <= execute_ctrl2_down_RS2_RFID_lane0;
      execute_ctrl3_up_RS2_PHYS_lane0 <= execute_ctrl2_down_RS2_PHYS_lane0;
      execute_ctrl3_up_RD_ENABLE_lane0 <= execute_ctrl2_down_RD_ENABLE_lane0;
      execute_ctrl3_up_RD_RFID_lane0 <= execute_ctrl2_down_RD_RFID_lane0;
      execute_ctrl3_up_RD_PHYS_lane0 <= execute_ctrl2_down_RD_PHYS_lane0;
      execute_ctrl3_up_LANE_AGE_lane0 <= execute_ctrl2_down_LANE_AGE_lane0;
      execute_ctrl3_up_COMPLETED_lane0 <= execute_ctrl2_down_COMPLETED_lane0;
      execute_ctrl3_up_Decode_UOP_lane1 <= execute_ctrl2_down_Decode_UOP_lane1;
      execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1 <= execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1;
      execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1 <= execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
      execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      execute_ctrl3_up_PC_lane1 <= execute_ctrl2_down_PC_lane1;
      execute_ctrl3_up_TRAP_lane1 <= execute_ctrl2_down_TRAP_lane1;
      execute_ctrl3_up_Decode_UOP_ID_lane1 <= execute_ctrl2_down_Decode_UOP_ID_lane1;
      execute_ctrl3_up_RS1_RFID_lane1 <= execute_ctrl2_down_RS1_RFID_lane1;
      execute_ctrl3_up_RS1_PHYS_lane1 <= execute_ctrl2_down_RS1_PHYS_lane1;
      execute_ctrl3_up_RS2_RFID_lane1 <= execute_ctrl2_down_RS2_RFID_lane1;
      execute_ctrl3_up_RS2_PHYS_lane1 <= execute_ctrl2_down_RS2_PHYS_lane1;
      execute_ctrl3_up_RD_ENABLE_lane1 <= execute_ctrl2_down_RD_ENABLE_lane1;
      execute_ctrl3_up_RD_RFID_lane1 <= execute_ctrl2_down_RD_RFID_lane1;
      execute_ctrl3_up_RD_PHYS_lane1 <= execute_ctrl2_down_RD_PHYS_lane1;
      execute_ctrl3_up_LANE_AGE_lane1 <= execute_ctrl2_down_LANE_AGE_lane1;
      execute_ctrl3_up_COMPLETED_lane1 <= execute_ctrl2_down_COMPLETED_lane1;
      execute_ctrl3_up_AguPlugin_SIZE_lane0 <= execute_ctrl2_down_AguPlugin_SIZE_lane0;
      execute_ctrl3_up_integer_RS1_lane0 <= execute_ctrl2_down_integer_RS1_lane0;
      execute_ctrl3_up_integer_RS2_lane0 <= execute_ctrl2_down_integer_RS2_lane0;
      execute_ctrl3_up_integer_RS1_lane1 <= execute_ctrl2_down_integer_RS1_lane1;
      execute_ctrl3_up_integer_RS2_lane1 <= execute_ctrl2_down_integer_RS2_lane1;
      execute_ctrl3_up_float_RS1_lane0 <= execute_ctrl2_down_float_RS1_lane0;
      execute_ctrl3_up_float_RS2_lane0 <= execute_ctrl2_down_float_RS2_lane0;
      execute_ctrl3_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl3_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl3_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0 <= execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0;
      execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl3_up_late0_BranchPlugin_SEL_lane0 <= execute_ctrl2_down_late0_BranchPlugin_SEL_lane0;
      execute_ctrl3_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl3_up_FpuCsrPlugin_DIRTY_lane0 <= execute_ctrl2_down_FpuCsrPlugin_DIRTY_lane0;
      execute_ctrl3_up_FpuClassPlugin_SEL_lane0 <= execute_ctrl2_down_FpuClassPlugin_SEL_lane0;
      execute_ctrl3_up_FpuCmpPlugin_SEL_FLOAT_lane0 <= execute_ctrl2_down_FpuCmpPlugin_SEL_FLOAT_lane0;
      execute_ctrl3_up_FpuCmpPlugin_SEL_CMP_lane0 <= execute_ctrl2_down_FpuCmpPlugin_SEL_CMP_lane0;
      execute_ctrl3_up_FpuF2iPlugin_SEL_lane0 <= execute_ctrl2_down_FpuF2iPlugin_SEL_lane0;
      execute_ctrl3_up_FpuMvPlugin_SEL_FLOAT_lane0 <= execute_ctrl2_down_FpuMvPlugin_SEL_FLOAT_lane0;
      execute_ctrl3_up_FpuMvPlugin_SEL_INT_lane0 <= execute_ctrl2_down_FpuMvPlugin_SEL_INT_lane0;
      execute_ctrl3_up_AguPlugin_SEL_lane0 <= execute_ctrl2_down_AguPlugin_SEL_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl3_up_FpuMulPlugin_SEL_lane0 <= execute_ctrl2_down_FpuMulPlugin_SEL_lane0;
      execute_ctrl3_up_FpuXxPlugin_SEL_lane0 <= execute_ctrl2_down_FpuXxPlugin_SEL_lane0;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl3_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl2_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl3_up_COMPLETION_AT_4_lane0 <= execute_ctrl2_down_COMPLETION_AT_4_lane0;
      execute_ctrl3_up_COMPLETION_AT_7_lane0 <= execute_ctrl2_down_COMPLETION_AT_7_lane0;
      execute_ctrl3_up_COMPLETION_AT_11_lane0 <= execute_ctrl2_down_COMPLETION_AT_11_lane0;
      execute_ctrl3_up_COMPLETION_AT_3_lane0 <= execute_ctrl2_down_COMPLETION_AT_3_lane0;
      execute_ctrl3_up_COMPLETION_AT_5_lane0 <= execute_ctrl2_down_COMPLETION_AT_5_lane0;
      execute_ctrl3_up_COMPLETION_AT_8_lane0 <= execute_ctrl2_down_COMPLETION_AT_8_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_3_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_3_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl3_up_SrcStageables_REVERT_lane0 <= execute_ctrl2_down_SrcStageables_REVERT_lane0;
      execute_ctrl3_up_SrcStageables_ZERO_lane0 <= execute_ctrl2_down_SrcStageables_ZERO_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl3_up_BYPASSED_AT_4_lane0 <= execute_ctrl2_down_BYPASSED_AT_4_lane0;
      execute_ctrl3_up_BYPASSED_AT_5_lane0 <= execute_ctrl2_down_BYPASSED_AT_5_lane0;
      execute_ctrl3_up_BYPASSED_AT_6_lane0 <= execute_ctrl2_down_BYPASSED_AT_6_lane0;
      execute_ctrl3_up_BYPASSED_AT_7_lane0 <= execute_ctrl2_down_BYPASSED_AT_7_lane0;
      execute_ctrl3_up_BYPASSED_AT_8_lane0 <= execute_ctrl2_down_BYPASSED_AT_8_lane0;
      execute_ctrl3_up_BYPASSED_AT_9_lane0 <= execute_ctrl2_down_BYPASSED_AT_9_lane0;
      execute_ctrl3_up_BYPASSED_AT_10_lane0 <= execute_ctrl2_down_BYPASSED_AT_10_lane0;
      execute_ctrl3_up_SrcStageables_UNSIGNED_lane0 <= execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
      execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0 <= execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
      execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0 <= execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
      execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl3_up_MulPlugin_HIGH_lane0 <= execute_ctrl2_down_MulPlugin_HIGH_lane0;
      execute_ctrl3_up_FpuUtils_FORMAT_lane0 <= execute_ctrl2_down_FpuUtils_FORMAT_lane0;
      execute_ctrl3_up_FpuCmpPlugin_FLOAT_OP_lane0 <= execute_ctrl2_down_FpuCmpPlugin_FLOAT_OP_lane0;
      execute_ctrl3_up_AguPlugin_LOAD_lane0 <= execute_ctrl2_down_AguPlugin_LOAD_lane0;
      execute_ctrl3_up_AguPlugin_STORE_lane0 <= execute_ctrl2_down_AguPlugin_STORE_lane0;
      execute_ctrl3_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl3_up_AguPlugin_FLOAT_lane0 <= execute_ctrl2_down_AguPlugin_FLOAT_lane0;
      execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl3_up_FpuMulPlugin_FMA_lane0 <= execute_ctrl2_down_FpuMulPlugin_FMA_lane0;
      execute_ctrl3_up_FpuMulPlugin_SUB1_lane0 <= execute_ctrl2_down_FpuMulPlugin_SUB1_lane0;
      execute_ctrl3_up_FpuMulPlugin_SUB2_lane0 <= execute_ctrl2_down_FpuMulPlugin_SUB2_lane0;
      execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0 <= execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
      execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0 <= execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
      execute_ctrl3_up_early1_BranchPlugin_SEL_lane1 <= execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
      execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1 <= execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1;
      execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1 <= execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1;
      execute_ctrl3_up_late1_BranchPlugin_SEL_lane1 <= execute_ctrl2_down_late1_BranchPlugin_SEL_lane1;
      execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      execute_ctrl3_up_COMPLETION_AT_4_lane1 <= execute_ctrl2_down_COMPLETION_AT_4_lane1;
      execute_ctrl3_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1 <= execute_ctrl2_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
      execute_ctrl3_up_SrcStageables_REVERT_lane1 <= execute_ctrl2_down_SrcStageables_REVERT_lane1;
      execute_ctrl3_up_SrcStageables_ZERO_lane1 <= execute_ctrl2_down_SrcStageables_ZERO_lane1;
      execute_ctrl3_up_SrcStageables_UNSIGNED_lane1 <= execute_ctrl2_down_SrcStageables_UNSIGNED_lane1;
      execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1 <= execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1;
      execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1 <= execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1;
      execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1 <= execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1;
      execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1 <= execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
      execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1 <= execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
      execute_ctrl3_up_COMMIT_lane0 <= execute_ctrl2_down_COMMIT_lane0;
      execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX <= execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
      execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF <= execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
      execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF <= execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
      execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ <= execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
      execute_ctrl3_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV <= execute_ctrl2_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
      execute_ctrl3_up_COMMIT_lane1 <= execute_ctrl2_down_COMMIT_lane1;
      execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0 <= execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
      execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_4_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_5_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_6_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_7_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_8_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_9_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_10_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_11_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_12_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_13_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_14_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_15_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
      execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0 <= execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
      execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 <= execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
      execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 <= execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
      execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 <= execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
      execute_ctrl3_up_FpuUtils_ROUNDING_lane0 <= execute_ctrl2_down_FpuUtils_ROUNDING_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_WB_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0;
      execute_ctrl3_up_LsuL1_MASK_lane0 <= execute_ctrl2_down_LsuL1_MASK_lane0;
      execute_ctrl3_up_LsuL1_SIZE_lane0 <= execute_ctrl2_down_LsuL1_SIZE_lane0;
      execute_ctrl3_up_LsuL1_LOAD_lane0 <= execute_ctrl2_down_LsuL1_LOAD_lane0;
      execute_ctrl3_up_LsuL1_ATOMIC_lane0 <= execute_ctrl2_down_LsuL1_ATOMIC_lane0;
      execute_ctrl3_up_LsuL1_STORE_lane0 <= execute_ctrl2_down_LsuL1_STORE_lane0;
      execute_ctrl3_up_LsuL1_CLEAN_lane0 <= execute_ctrl2_down_LsuL1_CLEAN_lane0;
      execute_ctrl3_up_LsuL1_INVALID_lane0 <= execute_ctrl2_down_LsuL1_INVALID_lane0;
      execute_ctrl3_up_LsuL1_PREFETCH_lane0 <= execute_ctrl2_down_LsuL1_PREFETCH_lane0;
      execute_ctrl3_up_LsuL1_FLUSH_lane0 <= execute_ctrl2_down_LsuL1_FLUSH_lane0;
      execute_ctrl3_up_Decode_STORE_ID_lane0 <= execute_ctrl2_down_Decode_STORE_ID_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl3_up_LsuPlugin_SB_PTR_lane0 <= execute_ctrl2_down_LsuPlugin_SB_PTR_lane0;
      execute_ctrl3_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0 <= execute_ctrl2_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
      execute_ctrl3_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0 <= execute_ctrl2_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
      execute_ctrl3_up_FpuUnpack_RS1_IS_SUBNORMAL_lane0 <= execute_ctrl2_down_FpuUnpack_RS1_IS_SUBNORMAL_lane0;
      execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mode <= execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mode;
      execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_quiet <= execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_quiet;
      execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_sign <= execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_sign;
      execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent <= _zz_execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_exponent;
      execute_ctrl3_up_FpuUnpack_RS1_RS_lane0_mantissa <= execute_ctrl2_down_FpuUnpack_RS1_RS_lane0_mantissa;
      execute_ctrl3_up_FpuUnpack_RS1_badBoxing_HIT_lane0 <= execute_ctrl2_down_FpuUnpack_RS1_badBoxing_HIT_lane0;
      execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mode <= execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mode;
      execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_quiet <= execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_quiet;
      execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_sign <= execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_sign;
      execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent <= _zz_execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_exponent;
      execute_ctrl3_up_FpuUnpack_RS2_RS_lane0_mantissa <= execute_ctrl2_down_FpuUnpack_RS2_RS_lane0_mantissa;
      execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mode <= execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mode;
      execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_quiet <= execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_quiet;
      execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_sign <= execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_sign;
      execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent <= _zz_execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_exponent;
      execute_ctrl3_up_FpuUnpack_RS3_RS_lane0_mantissa <= execute_ctrl2_down_FpuUnpack_RS3_RS_lane0_mantissa;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
      execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0 <= execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_MIN_MAX_RS2_lane0;
      execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0 <= execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_CMP_RESULT_lane0;
      execute_ctrl3_up_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0 <= execute_ctrl2_down_FpuCmpPlugin_logic_onCmp_SGNJ_RESULT_lane0;
      execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_f2iShift_lane0 <= execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_f2iShift_lane0;
      execute_ctrl3_up_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0 <= execute_ctrl2_down_FpuF2iPlugin_logic_onSetup_SHIFTED_PARTIAL_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 <= _zz_execute_ctrl3_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_SIGN_lane0 <= execute_ctrl2_down_FpuMulPlugin_logic_calc_SIGN_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 <= execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 <= execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 <= execute_ctrl2_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
      execute_ctrl3_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 <= execute_ctrl2_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
    end
    if(execute_ctrl3_down_isReady) begin
      execute_ctrl4_up_Decode_UOP_lane0 <= execute_ctrl3_down_Decode_UOP_lane0;
      execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0 <= execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_6_lane0;
      execute_ctrl4_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl3_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl4_up_PC_lane0 <= execute_ctrl3_down_PC_lane0;
      execute_ctrl4_up_TRAP_lane0 <= execute_ctrl3_down_TRAP_lane0;
      execute_ctrl4_up_Decode_UOP_ID_lane0 <= execute_ctrl3_down_Decode_UOP_ID_lane0;
      execute_ctrl4_up_RD_ENABLE_lane0 <= execute_ctrl3_down_RD_ENABLE_lane0;
      execute_ctrl4_up_RD_RFID_lane0 <= execute_ctrl3_down_RD_RFID_lane0;
      execute_ctrl4_up_RD_PHYS_lane0 <= execute_ctrl3_down_RD_PHYS_lane0;
      execute_ctrl4_up_LANE_AGE_lane0 <= execute_ctrl3_down_LANE_AGE_lane0;
      execute_ctrl4_up_COMPLETED_lane0 <= execute_ctrl3_down_COMPLETED_lane0;
      execute_ctrl4_up_Decode_UOP_lane1 <= execute_ctrl3_down_Decode_UOP_lane1;
      execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1 <= execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1;
      execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1 <= execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
      execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      execute_ctrl4_up_PC_lane1 <= execute_ctrl3_down_PC_lane1;
      execute_ctrl4_up_TRAP_lane1 <= execute_ctrl3_down_TRAP_lane1;
      execute_ctrl4_up_Decode_UOP_ID_lane1 <= execute_ctrl3_down_Decode_UOP_ID_lane1;
      execute_ctrl4_up_RD_ENABLE_lane1 <= execute_ctrl3_down_RD_ENABLE_lane1;
      execute_ctrl4_up_RD_RFID_lane1 <= execute_ctrl3_down_RD_RFID_lane1;
      execute_ctrl4_up_RD_PHYS_lane1 <= execute_ctrl3_down_RD_PHYS_lane1;
      execute_ctrl4_up_LANE_AGE_lane1 <= execute_ctrl3_down_LANE_AGE_lane1;
      execute_ctrl4_up_COMPLETED_lane1 <= execute_ctrl3_down_COMPLETED_lane1;
      execute_ctrl4_up_AguPlugin_SIZE_lane0 <= execute_ctrl3_down_AguPlugin_SIZE_lane0;
      execute_ctrl4_up_integer_RS1_lane0 <= execute_ctrl3_down_integer_RS1_lane0;
      execute_ctrl4_up_integer_RS2_lane0 <= execute_ctrl3_down_integer_RS2_lane0;
      execute_ctrl4_up_float_RS2_lane0 <= execute_ctrl3_down_float_RS2_lane0;
      execute_ctrl4_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl3_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl4_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0 <= execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0;
      execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl4_up_late0_BranchPlugin_SEL_lane0 <= execute_ctrl3_down_late0_BranchPlugin_SEL_lane0;
      execute_ctrl4_up_FpuCsrPlugin_DIRTY_lane0 <= execute_ctrl3_down_FpuCsrPlugin_DIRTY_lane0;
      execute_ctrl4_up_FpuF2iPlugin_SEL_lane0 <= execute_ctrl3_down_FpuF2iPlugin_SEL_lane0;
      execute_ctrl4_up_FpuMvPlugin_SEL_FLOAT_lane0 <= execute_ctrl3_down_FpuMvPlugin_SEL_FLOAT_lane0;
      execute_ctrl4_up_AguPlugin_SEL_lane0 <= execute_ctrl3_down_AguPlugin_SEL_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl4_up_FpuMulPlugin_SEL_lane0 <= execute_ctrl3_down_FpuMulPlugin_SEL_lane0;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl4_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl3_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl4_up_COMPLETION_AT_4_lane0 <= execute_ctrl3_down_COMPLETION_AT_4_lane0;
      execute_ctrl4_up_COMPLETION_AT_7_lane0 <= execute_ctrl3_down_COMPLETION_AT_7_lane0;
      execute_ctrl4_up_COMPLETION_AT_11_lane0 <= execute_ctrl3_down_COMPLETION_AT_11_lane0;
      execute_ctrl4_up_COMPLETION_AT_5_lane0 <= execute_ctrl3_down_COMPLETION_AT_5_lane0;
      execute_ctrl4_up_COMPLETION_AT_8_lane0 <= execute_ctrl3_down_COMPLETION_AT_8_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl4_up_SrcStageables_REVERT_lane0 <= execute_ctrl3_down_SrcStageables_REVERT_lane0;
      execute_ctrl4_up_SrcStageables_ZERO_lane0 <= execute_ctrl3_down_SrcStageables_ZERO_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl4_up_BYPASSED_AT_5_lane0 <= execute_ctrl3_down_BYPASSED_AT_5_lane0;
      execute_ctrl4_up_BYPASSED_AT_6_lane0 <= execute_ctrl3_down_BYPASSED_AT_6_lane0;
      execute_ctrl4_up_BYPASSED_AT_7_lane0 <= execute_ctrl3_down_BYPASSED_AT_7_lane0;
      execute_ctrl4_up_BYPASSED_AT_8_lane0 <= execute_ctrl3_down_BYPASSED_AT_8_lane0;
      execute_ctrl4_up_BYPASSED_AT_9_lane0 <= execute_ctrl3_down_BYPASSED_AT_9_lane0;
      execute_ctrl4_up_BYPASSED_AT_10_lane0 <= execute_ctrl3_down_BYPASSED_AT_10_lane0;
      execute_ctrl4_up_SrcStageables_UNSIGNED_lane0 <= execute_ctrl3_down_SrcStageables_UNSIGNED_lane0;
      execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0 <= execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0;
      execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0 <= execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0;
      execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl4_up_MulPlugin_HIGH_lane0 <= execute_ctrl3_down_MulPlugin_HIGH_lane0;
      execute_ctrl4_up_FpuUtils_FORMAT_lane0 <= execute_ctrl3_down_FpuUtils_FORMAT_lane0;
      execute_ctrl4_up_AguPlugin_LOAD_lane0 <= execute_ctrl3_down_AguPlugin_LOAD_lane0;
      execute_ctrl4_up_AguPlugin_STORE_lane0 <= execute_ctrl3_down_AguPlugin_STORE_lane0;
      execute_ctrl4_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl4_up_AguPlugin_FLOAT_lane0 <= execute_ctrl3_down_AguPlugin_FLOAT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl4_up_FpuMulPlugin_FMA_lane0 <= execute_ctrl3_down_FpuMulPlugin_FMA_lane0;
      execute_ctrl4_up_FpuMulPlugin_SUB1_lane0 <= execute_ctrl3_down_FpuMulPlugin_SUB1_lane0;
      execute_ctrl4_up_FpuMulPlugin_SUB2_lane0 <= execute_ctrl3_down_FpuMulPlugin_SUB2_lane0;
      execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl4_up_early1_BranchPlugin_SEL_lane1 <= execute_ctrl3_down_early1_BranchPlugin_SEL_lane1;
      execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1 <= execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1;
      execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1 <= execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1;
      execute_ctrl4_up_late1_BranchPlugin_SEL_lane1 <= execute_ctrl3_down_late1_BranchPlugin_SEL_lane1;
      execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      execute_ctrl4_up_COMPLETION_AT_4_lane1 <= execute_ctrl3_down_COMPLETION_AT_4_lane1;
      execute_ctrl4_up_lane1_logic_completions_onCtrl_1_ENABLE_lane1 <= execute_ctrl3_down_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
      execute_ctrl4_up_SrcStageables_REVERT_lane1 <= execute_ctrl3_down_SrcStageables_REVERT_lane1;
      execute_ctrl4_up_SrcStageables_ZERO_lane1 <= execute_ctrl3_down_SrcStageables_ZERO_lane1;
      execute_ctrl4_up_SrcStageables_UNSIGNED_lane1 <= execute_ctrl3_down_SrcStageables_UNSIGNED_lane1;
      execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1 <= execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1;
      execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1 <= execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1;
      execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1 <= execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1;
      execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      execute_ctrl4_up_COMMIT_lane0 <= execute_ctrl3_down_COMMIT_lane0;
      execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX <= execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NX;
      execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF <= execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_UF;
      execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF <= execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_OF;
      execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ <= execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_DZ;
      execute_ctrl4_up_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV <= execute_ctrl3_down_FpuFlagsWritebackPlugin_logic_FLAGS_lane0_NV;
      execute_ctrl4_up_COMMIT_lane1 <= execute_ctrl3_down_COMMIT_lane1;
      execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_4_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_4_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_5_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_5_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_6_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_6_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_7_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_7_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_8_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_8_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_9_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_9_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_10_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_10_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_11_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_11_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_12_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_12_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_13_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_13_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_14_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_14_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_15_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_15_lane0;
      execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 <= execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
      execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 <= execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
      execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 <= execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
      execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 <= execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
      execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 <= execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
      execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 <= execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
      execute_ctrl4_up_FpuUtils_ROUNDING_lane0 <= execute_ctrl3_down_FpuUtils_ROUNDING_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_WB_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_WB_lane0;
      execute_ctrl4_up_LsuL1_MASK_lane0 <= execute_ctrl3_down_LsuL1_MASK_lane0;
      execute_ctrl4_up_LsuL1_SIZE_lane0 <= execute_ctrl3_down_LsuL1_SIZE_lane0;
      execute_ctrl4_up_LsuL1_LOAD_lane0 <= execute_ctrl3_down_LsuL1_LOAD_lane0;
      execute_ctrl4_up_LsuL1_ATOMIC_lane0 <= execute_ctrl3_down_LsuL1_ATOMIC_lane0;
      execute_ctrl4_up_LsuL1_STORE_lane0 <= execute_ctrl3_down_LsuL1_STORE_lane0;
      execute_ctrl4_up_LsuL1_CLEAN_lane0 <= execute_ctrl3_down_LsuL1_CLEAN_lane0;
      execute_ctrl4_up_LsuL1_INVALID_lane0 <= execute_ctrl3_down_LsuL1_INVALID_lane0;
      execute_ctrl4_up_LsuL1_PREFETCH_lane0 <= execute_ctrl3_down_LsuL1_PREFETCH_lane0;
      execute_ctrl4_up_LsuL1_FLUSH_lane0 <= execute_ctrl3_down_LsuL1_FLUSH_lane0;
      execute_ctrl4_up_Decode_STORE_ID_lane0 <= execute_ctrl3_down_Decode_STORE_ID_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl4_up_LsuPlugin_SB_PTR_lane0 <= execute_ctrl3_down_LsuPlugin_SB_PTR_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onAddress0_SB_DATA_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onAddress0_SB_DATA_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onAddress0_STORE_BUFFER_EMPTY_lane0;
      execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mode <= execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mode;
      execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_quiet <= execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_quiet;
      execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_sign <= execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_sign;
      execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent <= _zz_execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_exponent;
      execute_ctrl4_up_FpuUnpack_RS1_RS_lane0_mantissa <= execute_ctrl3_down_FpuUnpack_RS1_RS_lane0_mantissa;
      execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mode <= execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mode;
      execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_quiet <= execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_quiet;
      execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_sign <= execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_sign;
      execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent <= _zz_execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_exponent;
      execute_ctrl4_up_FpuUnpack_RS2_RS_lane0_mantissa <= execute_ctrl3_down_FpuUnpack_RS2_RS_lane0_mantissa;
      execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mode <= execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mode;
      execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_quiet <= execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_quiet;
      execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_sign <= execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_sign;
      execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent <= _zz_execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_exponent;
      execute_ctrl4_up_FpuUnpack_RS3_RS_lane0_mantissa <= execute_ctrl3_down_FpuUnpack_RS3_RS_lane0_mantissa;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 <= _zz_execute_ctrl4_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_SIGN_lane0 <= execute_ctrl3_down_FpuMulPlugin_logic_calc_SIGN_lane0;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 <= execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 <= execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 <= execute_ctrl3_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
      execute_ctrl4_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 <= execute_ctrl3_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
      execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
      execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
      execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
      execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0 <= execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
      execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0 <= execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
      execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1 <= execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
      execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1 <= execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_2_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_2_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
      execute_ctrl4_up_MMU_TRANSLATED_lane0 <= execute_ctrl3_down_MMU_TRANSLATED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
      execute_ctrl4_up_MMU_ACCESS_FAULT_lane0 <= execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
      execute_ctrl4_up_MMU_REFILL_lane0 <= execute_ctrl3_down_MMU_REFILL_lane0;
      execute_ctrl4_up_MMU_HAZARD_lane0 <= execute_ctrl3_down_MMU_HAZARD_lane0;
      execute_ctrl4_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl3_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl4_up_FpuF2iPlugin_logic_onShift_SHIFTED_lane0 <= execute_ctrl3_down_FpuF2iPlugin_logic_onShift_SHIFTED_lane0;
      execute_ctrl4_up_FpuF2iPlugin_logic_onShift_resign_lane0 <= execute_ctrl3_down_FpuF2iPlugin_logic_onShift_resign_lane0;
      execute_ctrl4_up_FpuF2iPlugin_logic_onShift_increment_lane0 <= execute_ctrl3_down_FpuF2iPlugin_logic_onShift_increment_lane0;
      execute_ctrl4_up_FpuF2iPlugin_logic_onShift_incrementPatched_lane0 <= execute_ctrl3_down_FpuF2iPlugin_logic_onShift_incrementPatched_lane0;
      execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0 <= execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
    end
    if(execute_ctrl4_down_isReady) begin
      execute_ctrl5_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl4_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl5_up_TRAP_lane0 <= execute_ctrl4_down_TRAP_lane0;
      execute_ctrl5_up_Decode_UOP_ID_lane0 <= execute_ctrl4_down_Decode_UOP_ID_lane0;
      execute_ctrl5_up_RD_ENABLE_lane0 <= execute_ctrl4_down_RD_ENABLE_lane0;
      execute_ctrl5_up_RD_RFID_lane0 <= execute_ctrl4_down_RD_RFID_lane0;
      execute_ctrl5_up_RD_PHYS_lane0 <= execute_ctrl4_down_RD_PHYS_lane0;
      execute_ctrl5_up_LANE_AGE_lane0 <= execute_ctrl4_down_LANE_AGE_lane0;
      execute_ctrl5_up_COMPLETED_lane0 <= execute_ctrl4_down_COMPLETED_lane0;
      execute_ctrl5_up_RD_ENABLE_lane1 <= execute_ctrl4_down_RD_ENABLE_lane1;
      execute_ctrl5_up_RD_RFID_lane1 <= execute_ctrl4_down_RD_RFID_lane1;
      execute_ctrl5_up_RD_PHYS_lane1 <= execute_ctrl4_down_RD_PHYS_lane1;
      execute_ctrl5_up_LANE_AGE_lane1 <= execute_ctrl4_down_LANE_AGE_lane1;
      execute_ctrl5_up_FpuMulPlugin_SEL_lane0 <= execute_ctrl4_down_FpuMulPlugin_SEL_lane0;
      execute_ctrl5_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl4_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl5_up_COMPLETION_AT_7_lane0 <= execute_ctrl4_down_COMPLETION_AT_7_lane0;
      execute_ctrl5_up_COMPLETION_AT_11_lane0 <= execute_ctrl4_down_COMPLETION_AT_11_lane0;
      execute_ctrl5_up_COMPLETION_AT_5_lane0 <= execute_ctrl4_down_COMPLETION_AT_5_lane0;
      execute_ctrl5_up_COMPLETION_AT_8_lane0 <= execute_ctrl4_down_COMPLETION_AT_8_lane0;
      execute_ctrl5_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl4_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl5_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl5_up_lane0_logic_completions_onCtrl_4_ENABLE_lane0 <= execute_ctrl4_down_lane0_logic_completions_onCtrl_4_ENABLE_lane0;
      execute_ctrl5_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl4_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl5_up_BYPASSED_AT_6_lane0 <= execute_ctrl4_down_BYPASSED_AT_6_lane0;
      execute_ctrl5_up_BYPASSED_AT_7_lane0 <= execute_ctrl4_down_BYPASSED_AT_7_lane0;
      execute_ctrl5_up_BYPASSED_AT_8_lane0 <= execute_ctrl4_down_BYPASSED_AT_8_lane0;
      execute_ctrl5_up_BYPASSED_AT_9_lane0 <= execute_ctrl4_down_BYPASSED_AT_9_lane0;
      execute_ctrl5_up_BYPASSED_AT_10_lane0 <= execute_ctrl4_down_BYPASSED_AT_10_lane0;
      execute_ctrl5_up_FpuUtils_FORMAT_lane0 <= execute_ctrl4_down_FpuUtils_FORMAT_lane0;
      execute_ctrl5_up_FpuMulPlugin_FMA_lane0 <= execute_ctrl4_down_FpuMulPlugin_FMA_lane0;
      execute_ctrl5_up_FpuMulPlugin_SUB1_lane0 <= execute_ctrl4_down_FpuMulPlugin_SUB1_lane0;
      execute_ctrl5_up_FpuMulPlugin_SUB2_lane0 <= execute_ctrl4_down_FpuMulPlugin_SUB2_lane0;
      execute_ctrl5_up_COMMIT_lane0 <= execute_ctrl4_down_COMMIT_lane0;
      execute_ctrl5_up_COMMIT_lane1 <= execute_ctrl4_down_COMMIT_lane1;
      execute_ctrl5_up_FpuUtils_ROUNDING_lane0 <= execute_ctrl4_down_FpuUtils_ROUNDING_lane0;
      execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mode <= execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mode;
      execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_quiet <= execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_quiet;
      execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_sign <= execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_sign;
      execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent <= _zz_execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_exponent;
      execute_ctrl5_up_FpuUnpack_RS1_RS_lane0_mantissa <= execute_ctrl4_down_FpuUnpack_RS1_RS_lane0_mantissa;
      execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mode <= execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mode;
      execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_quiet <= execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_quiet;
      execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_sign <= execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_sign;
      execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent <= _zz_execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_exponent;
      execute_ctrl5_up_FpuUnpack_RS2_RS_lane0_mantissa <= execute_ctrl4_down_FpuUnpack_RS2_RS_lane0_mantissa;
      execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mode <= execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mode;
      execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_quiet <= execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_quiet;
      execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_sign <= execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_sign;
      execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent <= _zz_execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_exponent;
      execute_ctrl5_up_FpuUnpack_RS3_RS_lane0_mantissa <= execute_ctrl4_down_FpuUnpack_RS3_RS_lane0_mantissa;
      execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0 <= _zz_execute_ctrl5_up_FpuMulPlugin_logic_calc_EXP_ADD_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_SIGN_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_calc_SIGN_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_ZERO_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_OVERFLOW_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_calc_INFINITY_NAN_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_calc_FORCE_NAN_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_calc_FORCE_NAN_lane0;
      execute_ctrl5_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl4_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl5_up_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0 <= execute_ctrl4_down_FpuMulPlugin_logic_mulRsp_MUL_RESULT_lane0;
    end
    if(execute_ctrl5_down_isReady) begin
      execute_ctrl6_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl5_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl6_up_TRAP_lane0 <= execute_ctrl5_down_TRAP_lane0;
      execute_ctrl6_up_Decode_UOP_ID_lane0 <= execute_ctrl5_down_Decode_UOP_ID_lane0;
      execute_ctrl6_up_RD_ENABLE_lane0 <= execute_ctrl5_down_RD_ENABLE_lane0;
      execute_ctrl6_up_RD_RFID_lane0 <= execute_ctrl5_down_RD_RFID_lane0;
      execute_ctrl6_up_RD_PHYS_lane0 <= execute_ctrl5_down_RD_PHYS_lane0;
      execute_ctrl6_up_LANE_AGE_lane0 <= execute_ctrl5_down_LANE_AGE_lane0;
      execute_ctrl6_up_COMPLETED_lane0 <= execute_ctrl5_down_COMPLETED_lane0;
      execute_ctrl6_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl5_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl6_up_COMPLETION_AT_7_lane0 <= execute_ctrl5_down_COMPLETION_AT_7_lane0;
      execute_ctrl6_up_COMPLETION_AT_11_lane0 <= execute_ctrl5_down_COMPLETION_AT_11_lane0;
      execute_ctrl6_up_COMPLETION_AT_8_lane0 <= execute_ctrl5_down_COMPLETION_AT_8_lane0;
      execute_ctrl6_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl5_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl6_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl5_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl6_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl5_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl6_up_BYPASSED_AT_7_lane0 <= execute_ctrl5_down_BYPASSED_AT_7_lane0;
      execute_ctrl6_up_BYPASSED_AT_8_lane0 <= execute_ctrl5_down_BYPASSED_AT_8_lane0;
      execute_ctrl6_up_BYPASSED_AT_9_lane0 <= execute_ctrl5_down_BYPASSED_AT_9_lane0;
      execute_ctrl6_up_BYPASSED_AT_10_lane0 <= execute_ctrl5_down_BYPASSED_AT_10_lane0;
      execute_ctrl6_up_COMMIT_lane0 <= execute_ctrl5_down_COMMIT_lane0;
      execute_ctrl6_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl5_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl6_down_isReady) begin
      execute_ctrl7_up_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0 <= execute_ctrl6_down_FpuPackerPlugin_RESERVED_ON_early0_AT_9_lane0;
      execute_ctrl7_up_TRAP_lane0 <= execute_ctrl6_down_TRAP_lane0;
      execute_ctrl7_up_Decode_UOP_ID_lane0 <= execute_ctrl6_down_Decode_UOP_ID_lane0;
      execute_ctrl7_up_RD_ENABLE_lane0 <= execute_ctrl6_down_RD_ENABLE_lane0;
      execute_ctrl7_up_RD_RFID_lane0 <= execute_ctrl6_down_RD_RFID_lane0;
      execute_ctrl7_up_RD_PHYS_lane0 <= execute_ctrl6_down_RD_PHYS_lane0;
      execute_ctrl7_up_LANE_AGE_lane0 <= execute_ctrl6_down_LANE_AGE_lane0;
      execute_ctrl7_up_COMPLETED_lane0 <= execute_ctrl6_down_COMPLETED_lane0;
      execute_ctrl7_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl6_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl7_up_COMPLETION_AT_7_lane0 <= execute_ctrl6_down_COMPLETION_AT_7_lane0;
      execute_ctrl7_up_COMPLETION_AT_11_lane0 <= execute_ctrl6_down_COMPLETION_AT_11_lane0;
      execute_ctrl7_up_COMPLETION_AT_8_lane0 <= execute_ctrl6_down_COMPLETION_AT_8_lane0;
      execute_ctrl7_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl6_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl7_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl6_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl7_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl6_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl7_up_BYPASSED_AT_8_lane0 <= execute_ctrl6_down_BYPASSED_AT_8_lane0;
      execute_ctrl7_up_BYPASSED_AT_9_lane0 <= execute_ctrl6_down_BYPASSED_AT_9_lane0;
      execute_ctrl7_up_BYPASSED_AT_10_lane0 <= execute_ctrl6_down_BYPASSED_AT_10_lane0;
      execute_ctrl7_up_COMMIT_lane0 <= execute_ctrl6_down_COMMIT_lane0;
      execute_ctrl7_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl6_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl7_down_isReady) begin
      execute_ctrl8_up_TRAP_lane0 <= execute_ctrl7_down_TRAP_lane0;
      execute_ctrl8_up_Decode_UOP_ID_lane0 <= execute_ctrl7_down_Decode_UOP_ID_lane0;
      execute_ctrl8_up_RD_ENABLE_lane0 <= execute_ctrl7_down_RD_ENABLE_lane0;
      execute_ctrl8_up_RD_RFID_lane0 <= execute_ctrl7_down_RD_RFID_lane0;
      execute_ctrl8_up_RD_PHYS_lane0 <= execute_ctrl7_down_RD_PHYS_lane0;
      execute_ctrl8_up_LANE_AGE_lane0 <= execute_ctrl7_down_LANE_AGE_lane0;
      execute_ctrl8_up_COMPLETED_lane0 <= execute_ctrl7_down_COMPLETED_lane0;
      execute_ctrl8_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl7_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl8_up_COMPLETION_AT_11_lane0 <= execute_ctrl7_down_COMPLETION_AT_11_lane0;
      execute_ctrl8_up_COMPLETION_AT_8_lane0 <= execute_ctrl7_down_COMPLETION_AT_8_lane0;
      execute_ctrl8_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl7_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl8_up_lane0_logic_completions_onCtrl_5_ENABLE_lane0 <= execute_ctrl7_down_lane0_logic_completions_onCtrl_5_ENABLE_lane0;
      execute_ctrl8_up_BYPASSED_AT_9_lane0 <= execute_ctrl7_down_BYPASSED_AT_9_lane0;
      execute_ctrl8_up_BYPASSED_AT_10_lane0 <= execute_ctrl7_down_BYPASSED_AT_10_lane0;
      execute_ctrl8_up_COMMIT_lane0 <= execute_ctrl7_down_COMMIT_lane0;
      execute_ctrl8_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl7_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl8_down_isReady) begin
      execute_ctrl9_up_TRAP_lane0 <= execute_ctrl8_down_TRAP_lane0;
      execute_ctrl9_up_Decode_UOP_ID_lane0 <= execute_ctrl8_down_Decode_UOP_ID_lane0;
      execute_ctrl9_up_RD_ENABLE_lane0 <= execute_ctrl8_down_RD_ENABLE_lane0;
      execute_ctrl9_up_RD_RFID_lane0 <= execute_ctrl8_down_RD_RFID_lane0;
      execute_ctrl9_up_RD_PHYS_lane0 <= execute_ctrl8_down_RD_PHYS_lane0;
      execute_ctrl9_up_LANE_AGE_lane0 <= execute_ctrl8_down_LANE_AGE_lane0;
      execute_ctrl9_up_COMPLETED_lane0 <= execute_ctrl8_down_COMPLETED_lane0;
      execute_ctrl9_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl8_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl9_up_COMPLETION_AT_11_lane0 <= execute_ctrl8_down_COMPLETION_AT_11_lane0;
      execute_ctrl9_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl8_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl9_up_BYPASSED_AT_10_lane0 <= execute_ctrl8_down_BYPASSED_AT_10_lane0;
      execute_ctrl9_up_COMMIT_lane0 <= execute_ctrl8_down_COMMIT_lane0;
      execute_ctrl9_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl8_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl9_down_isReady) begin
      execute_ctrl10_up_TRAP_lane0 <= execute_ctrl9_down_TRAP_lane0;
      execute_ctrl10_up_Decode_UOP_ID_lane0 <= execute_ctrl9_down_Decode_UOP_ID_lane0;
      execute_ctrl10_up_RD_ENABLE_lane0 <= execute_ctrl9_down_RD_ENABLE_lane0;
      execute_ctrl10_up_RD_RFID_lane0 <= execute_ctrl9_down_RD_RFID_lane0;
      execute_ctrl10_up_RD_PHYS_lane0 <= execute_ctrl9_down_RD_PHYS_lane0;
      execute_ctrl10_up_LANE_AGE_lane0 <= execute_ctrl9_down_LANE_AGE_lane0;
      execute_ctrl10_up_COMPLETED_lane0 <= execute_ctrl9_down_COMPLETED_lane0;
      execute_ctrl10_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl9_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl10_up_COMPLETION_AT_11_lane0 <= execute_ctrl9_down_COMPLETION_AT_11_lane0;
      execute_ctrl10_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl9_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl10_up_COMMIT_lane0 <= execute_ctrl9_down_COMMIT_lane0;
      execute_ctrl10_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl9_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl10_down_isReady) begin
      execute_ctrl11_up_TRAP_lane0 <= execute_ctrl10_down_TRAP_lane0;
      execute_ctrl11_up_Decode_UOP_ID_lane0 <= execute_ctrl10_down_Decode_UOP_ID_lane0;
      execute_ctrl11_up_RD_ENABLE_lane0 <= execute_ctrl10_down_RD_ENABLE_lane0;
      execute_ctrl11_up_RD_RFID_lane0 <= execute_ctrl10_down_RD_RFID_lane0;
      execute_ctrl11_up_RD_PHYS_lane0 <= execute_ctrl10_down_RD_PHYS_lane0;
      execute_ctrl11_up_LANE_AGE_lane0 <= execute_ctrl10_down_LANE_AGE_lane0;
      execute_ctrl11_up_COMPLETED_lane0 <= execute_ctrl10_down_COMPLETED_lane0;
      execute_ctrl11_up_lane0_float_WriteBackPlugin_SEL_lane0 <= execute_ctrl10_down_lane0_float_WriteBackPlugin_SEL_lane0;
      execute_ctrl11_up_COMPLETION_AT_11_lane0 <= execute_ctrl10_down_COMPLETION_AT_11_lane0;
      execute_ctrl11_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl10_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl11_up_COMMIT_lane0 <= execute_ctrl10_down_COMMIT_lane0;
      execute_ctrl11_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl10_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    if(execute_ctrl11_down_isReady) begin
      execute_ctrl12_up_RD_ENABLE_lane0 <= execute_ctrl11_down_RD_ENABLE_lane0;
      execute_ctrl12_up_RD_RFID_lane0 <= execute_ctrl11_down_RD_RFID_lane0;
      execute_ctrl12_up_RD_PHYS_lane0 <= execute_ctrl11_down_RD_PHYS_lane0;
      execute_ctrl12_up_LANE_AGE_lane0 <= execute_ctrl11_down_LANE_AGE_lane0;
      execute_ctrl12_up_lane0_float_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl11_down_lane0_float_WriteBackPlugin_logic_DATA_lane0;
    end
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_SB_DRAIN : begin
      end
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l363) begin
          LsuPlugin_logic_flusher_waiter <= LsuL1_WRITEBACK_BUSY;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        LsuPlugin_logic_flusher_waiter <= (LsuPlugin_logic_flusher_waiter & LsuL1_WRITEBACK_BUSY);
      end
      default : begin
        LsuPlugin_logic_flusher_cmdCounter <= 7'h0;
      end
    endcase
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_COMPUTE : begin
        TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg <= TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_interface_aluInput <= CsrAccessPlugin_bus_read_toWriteBits;
        CsrAccessPlugin_logic_fsm_interface_csrValue <= CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        REG_CSR_2047 <= COMB_CSR_2047;
        REG_CSR_1952 <= COMB_CSR_1952;
        REG_CSR_1953 <= COMB_CSR_1953;
        REG_CSR_1954 <= COMB_CSR_1954;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_3 <= COMB_CSR_3;
        REG_CSR_2 <= COMB_CSR_2;
        REG_CSR_1 <= COMB_CSR_1;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
        REG_CSR_FpuCsrPlugin_logic_csrDirty <= COMB_CSR_FpuCsrPlugin_logic_csrDirty;
        REG_CSR_CsrRamPlugin_csrMapper_selFilter <= COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
        REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter <= COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
      end
    endcase
  end


endmodule

module RegFileMem_1 (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_address,
  input  wire [63:0]   io_writes_0_data,
  input  wire [15:0]   io_writes_0_uopId,
  input  wire          io_reads_0_valid,
  input  wire [4:0]    io_reads_0_address,
  output wire [63:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [4:0]    io_reads_1_address,
  output wire [63:0]   io_reads_1_data,
  input  wire          io_reads_2_valid,
  input  wire [4:0]    io_reads_2_address,
  output wire [63:0]   io_reads_2_data,
  input  wire          clk,
  input  wire          reset
);

  reg        [63:0]   asMem_ram_spinal_port1;
  reg        [63:0]   asMem_ram_spinal_port2;
  reg        [63:0]   asMem_ram_spinal_port3;
  reg                 _zz_1;
  wire                conv_writes_0_valid;
  wire       [4:0]    conv_writes_0_payload_address;
  wire       [63:0]   conv_writes_0_payload_data;
  wire                conv_read_0_cmd_valid;
  wire       [4:0]    conv_read_0_cmd_payload;
  wire       [63:0]   conv_read_0_rsp;
  wire                conv_read_1_cmd_valid;
  wire       [4:0]    conv_read_1_cmd_payload;
  wire       [63:0]   conv_read_1_rsp;
  wire                conv_read_2_cmd_valid;
  wire       [4:0]    conv_read_2_cmd_payload;
  wire       [63:0]   conv_read_2_rsp;
  wire                asMem_writes_0_port_valid;
  wire       [4:0]    asMem_writes_0_port_payload_address;
  wire       [63:0]   asMem_writes_0_port_payload_data;
  wire                asMem_reads_0_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_0_sync_port_cmd_payload;
  wire       [63:0]   asMem_reads_0_sync_port_rsp;
  wire                asMem_reads_1_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_1_sync_port_cmd_payload;
  wire       [63:0]   asMem_reads_1_sync_port_rsp;
  wire                asMem_reads_2_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_2_sync_port_cmd_payload;
  wire       [63:0]   asMem_reads_2_sync_port_rsp;
  reg [63:0] asMem_ram [0:31] /* verilator public */ ;

  always @(posedge clk) begin
    if(_zz_1) begin
      asMem_ram[asMem_writes_0_port_payload_address] <= asMem_writes_0_port_payload_data;
    end
  end

  always @(posedge clk) begin
    if(asMem_reads_0_sync_port_cmd_valid) begin
      asMem_ram_spinal_port1 <= asMem_ram[asMem_reads_0_sync_port_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(asMem_reads_1_sync_port_cmd_valid) begin
      asMem_ram_spinal_port2 <= asMem_ram[asMem_reads_1_sync_port_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(asMem_reads_2_sync_port_cmd_valid) begin
      asMem_ram_spinal_port3 <= asMem_ram[asMem_reads_2_sync_port_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(asMem_writes_0_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign conv_writes_0_valid = io_writes_0_valid;
  assign conv_writes_0_payload_address = io_writes_0_address;
  assign conv_writes_0_payload_data = io_writes_0_data;
  assign conv_read_0_cmd_valid = io_reads_0_valid;
  assign conv_read_0_cmd_payload = io_reads_0_address;
  assign io_reads_0_data = conv_read_0_rsp;
  assign conv_read_1_cmd_valid = io_reads_1_valid;
  assign conv_read_1_cmd_payload = io_reads_1_address;
  assign io_reads_1_data = conv_read_1_rsp;
  assign conv_read_2_cmd_valid = io_reads_2_valid;
  assign conv_read_2_cmd_payload = io_reads_2_address;
  assign io_reads_2_data = conv_read_2_rsp;
  assign asMem_writes_0_port_valid = conv_writes_0_valid;
  assign asMem_writes_0_port_payload_address = conv_writes_0_payload_address;
  assign asMem_writes_0_port_payload_data = conv_writes_0_payload_data;
  assign asMem_reads_0_sync_port_rsp = asMem_ram_spinal_port1;
  assign asMem_reads_0_sync_port_cmd_valid = conv_read_0_cmd_valid;
  assign asMem_reads_0_sync_port_cmd_payload = conv_read_0_cmd_payload;
  assign conv_read_0_rsp = asMem_reads_0_sync_port_rsp;
  assign asMem_reads_1_sync_port_rsp = asMem_ram_spinal_port2;
  assign asMem_reads_1_sync_port_cmd_valid = conv_read_1_cmd_valid;
  assign asMem_reads_1_sync_port_cmd_payload = conv_read_1_cmd_payload;
  assign conv_read_1_rsp = asMem_reads_1_sync_port_rsp;
  assign asMem_reads_2_sync_port_rsp = asMem_ram_spinal_port3;
  assign asMem_reads_2_sync_port_cmd_valid = conv_read_2_cmd_valid;
  assign asMem_reads_2_sync_port_cmd_payload = conv_read_2_cmd_payload;
  assign conv_read_2_rsp = asMem_reads_2_sync_port_rsp;

endmodule

module RegFileMem (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_address,
  input  wire [31:0]   io_writes_0_data,
  input  wire [15:0]   io_writes_0_uopId,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_address,
  input  wire [31:0]   io_writes_1_data,
  input  wire [15:0]   io_writes_1_uopId,
  input  wire          io_reads_0_valid,
  input  wire [4:0]    io_reads_0_address,
  output wire [31:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [4:0]    io_reads_1_address,
  output wire [31:0]   io_reads_1_data,
  input  wire          io_reads_2_valid,
  input  wire [4:0]    io_reads_2_address,
  output wire [31:0]   io_reads_2_data,
  input  wire          io_reads_3_valid,
  input  wire [4:0]    io_reads_3_address,
  output wire [31:0]   io_reads_3_data,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   ramSyncMwMux_1_io_read_0_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_1_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_2_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_3_rsp;
  wire                conv_writes_0_valid;
  wire       [4:0]    conv_writes_0_payload_address;
  wire       [31:0]   conv_writes_0_payload_data;
  wire                conv_writes_1_valid;
  wire       [4:0]    conv_writes_1_payload_address;
  wire       [31:0]   conv_writes_1_payload_data;
  wire                conv_read_0_cmd_valid;
  wire       [4:0]    conv_read_0_cmd_payload;
  wire       [31:0]   conv_read_0_rsp;
  wire                conv_read_1_cmd_valid;
  wire       [4:0]    conv_read_1_cmd_payload;
  wire       [31:0]   conv_read_1_rsp;
  wire                conv_read_2_cmd_valid;
  wire       [4:0]    conv_read_2_cmd_payload;
  wire       [31:0]   conv_read_2_rsp;
  wire                conv_read_3_cmd_valid;
  wire       [4:0]    conv_read_3_cmd_payload;
  wire       [31:0]   conv_read_3_rsp;

  RamSyncMwMux ramSyncMwMux_1 (
    .io_writes_0_valid           (conv_writes_0_valid               ), //i
    .io_writes_0_payload_address (conv_writes_0_payload_address[4:0]), //i
    .io_writes_0_payload_data    (conv_writes_0_payload_data[31:0]  ), //i
    .io_writes_1_valid           (conv_writes_1_valid               ), //i
    .io_writes_1_payload_address (conv_writes_1_payload_address[4:0]), //i
    .io_writes_1_payload_data    (conv_writes_1_payload_data[31:0]  ), //i
    .io_read_0_cmd_valid         (conv_read_0_cmd_valid             ), //i
    .io_read_0_cmd_payload       (conv_read_0_cmd_payload[4:0]      ), //i
    .io_read_0_rsp               (ramSyncMwMux_1_io_read_0_rsp[31:0]), //o
    .io_read_1_cmd_valid         (conv_read_1_cmd_valid             ), //i
    .io_read_1_cmd_payload       (conv_read_1_cmd_payload[4:0]      ), //i
    .io_read_1_rsp               (ramSyncMwMux_1_io_read_1_rsp[31:0]), //o
    .io_read_2_cmd_valid         (conv_read_2_cmd_valid             ), //i
    .io_read_2_cmd_payload       (conv_read_2_cmd_payload[4:0]      ), //i
    .io_read_2_rsp               (ramSyncMwMux_1_io_read_2_rsp[31:0]), //o
    .io_read_3_cmd_valid         (conv_read_3_cmd_valid             ), //i
    .io_read_3_cmd_payload       (conv_read_3_cmd_payload[4:0]      ), //i
    .io_read_3_rsp               (ramSyncMwMux_1_io_read_3_rsp[31:0]), //o
    .clk                         (clk                               ), //i
    .reset                       (reset                             )  //i
  );
  assign conv_writes_0_valid = io_writes_0_valid;
  assign conv_writes_0_payload_address = io_writes_0_address;
  assign conv_writes_0_payload_data = io_writes_0_data;
  assign conv_writes_1_valid = io_writes_1_valid;
  assign conv_writes_1_payload_address = io_writes_1_address;
  assign conv_writes_1_payload_data = io_writes_1_data;
  assign conv_read_0_cmd_valid = io_reads_0_valid;
  assign conv_read_0_cmd_payload = io_reads_0_address;
  assign io_reads_0_data = conv_read_0_rsp;
  assign conv_read_1_cmd_valid = io_reads_1_valid;
  assign conv_read_1_cmd_payload = io_reads_1_address;
  assign io_reads_1_data = conv_read_1_rsp;
  assign conv_read_2_cmd_valid = io_reads_2_valid;
  assign conv_read_2_cmd_payload = io_reads_2_address;
  assign io_reads_2_data = conv_read_2_rsp;
  assign conv_read_3_cmd_valid = io_reads_3_valid;
  assign conv_read_3_cmd_payload = io_reads_3_address;
  assign io_reads_3_data = conv_read_3_rsp;
  assign conv_read_0_rsp = ramSyncMwMux_1_io_read_0_rsp;
  assign conv_read_1_rsp = ramSyncMwMux_1_io_read_1_rsp;
  assign conv_read_2_rsp = ramSyncMwMux_1_io_read_2_rsp;
  assign conv_read_3_rsp = ramSyncMwMux_1_io_read_3_rsp;

endmodule

module FpuSqrt (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [53:0]   io_input_payload_a,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [52:0]   io_output_payload_result,
  output wire [56:0]   io_output_payload_remain,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);

  wire       [56:0]   _zz_t;
  wire       [54:0]   _zz_t_1;
  wire       [53:0]   _zz_q;
  wire       [58:0]   _zz_a_1;
  wire       [1:0]    _zz_a_2;
  reg        [5:0]    counter;
  reg                 busy;
  wire                io_output_fire;
  reg                 done;
  wire                when_FpuSqrt_l36;
  reg        [56:0]   a;
  reg        [51:0]   x;
  reg        [52:0]   q;
  wire       [56:0]   t;
  wire                when_FpuSqrt_l49;
  reg        [56:0]   _zz_a;
  wire                when_FpuSqrt_l52;
  wire                when_FpuSqrt_l60;

  assign _zz_t_1 = {q,2'b01};
  assign _zz_t = {2'd0, _zz_t_1};
  assign _zz_q = {q,(! t[56])};
  assign _zz_a_1 = {_zz_a,x[51 : 50]};
  assign _zz_a_2 = io_input_payload_a[53 : 52];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_FpuSqrt_l36 = (busy && (counter == 6'h35));
  assign t = (a - _zz_t);
  assign io_output_valid = done;
  assign io_output_payload_result = q;
  assign io_output_payload_remain = a;
  assign io_input_ready = (! busy);
  assign when_FpuSqrt_l49 = (! done);
  always @(*) begin
    _zz_a = a;
    if(when_FpuSqrt_l52) begin
      _zz_a = t;
    end
  end

  assign when_FpuSqrt_l52 = (! t[56]);
  assign when_FpuSqrt_l60 = (! busy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      busy <= 1'b0;
      done <= 1'b0;
    end else begin
      if(io_output_fire) begin
        busy <= 1'b0;
      end
      if(when_FpuSqrt_l36) begin
        done <= 1'b1;
      end
      if(io_output_fire) begin
        done <= 1'b0;
      end
      if(when_FpuSqrt_l60) begin
        if(io_input_valid) begin
          busy <= 1'b1;
        end
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_FpuSqrt_l49) begin
      counter <= (counter + 6'h01);
      q <= _zz_q[52:0];
      a <= _zz_a_1[56:0];
      x <= (x <<< 2);
    end
    if(when_FpuSqrt_l60) begin
      q <= 53'h0;
      a <= {55'd0, _zz_a_2};
      x <= io_input_payload_a[51:0];
      counter <= 6'h0;
    end
  end


endmodule

module StreamArbiter_4 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_pcOnLastSlice,
  input  wire [31:0]   io_inputs_0_payload_pcTarget,
  input  wire          io_inputs_0_payload_taken,
  input  wire          io_inputs_0_payload_isBranch,
  input  wire          io_inputs_0_payload_isPush,
  input  wire          io_inputs_0_payload_isPop,
  input  wire          io_inputs_0_payload_wasWrong,
  input  wire          io_inputs_0_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_0_payload_history,
  input  wire [15:0]   io_inputs_0_payload_uopId,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [31:0]   io_inputs_1_payload_pcOnLastSlice,
  input  wire [31:0]   io_inputs_1_payload_pcTarget,
  input  wire          io_inputs_1_payload_taken,
  input  wire          io_inputs_1_payload_isBranch,
  input  wire          io_inputs_1_payload_isPush,
  input  wire          io_inputs_1_payload_isPop,
  input  wire          io_inputs_1_payload_wasWrong,
  input  wire          io_inputs_1_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_1_payload_history,
  input  wire [15:0]   io_inputs_1_payload_uopId,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_pcOnLastSlice,
  output wire [31:0]   io_output_payload_pcTarget,
  output wire          io_output_payload_taken,
  output wire          io_output_payload_isBranch,
  output wire          io_output_payload_isPush,
  output wire          io_output_payload_isPop,
  output wire          io_output_payload_wasWrong,
  output wire          io_output_payload_badPredictedTarget,
  output wire [11:0]   io_output_payload_history,
  output wire [15:0]   io_output_payload_uopId,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_pcOnLastSlice = (maskRouted_0 ? io_inputs_0_payload_pcOnLastSlice : io_inputs_1_payload_pcOnLastSlice);
  assign io_output_payload_pcTarget = (maskRouted_0 ? io_inputs_0_payload_pcTarget : io_inputs_1_payload_pcTarget);
  assign io_output_payload_taken = (maskRouted_0 ? io_inputs_0_payload_taken : io_inputs_1_payload_taken);
  assign io_output_payload_isBranch = (maskRouted_0 ? io_inputs_0_payload_isBranch : io_inputs_1_payload_isBranch);
  assign io_output_payload_isPush = (maskRouted_0 ? io_inputs_0_payload_isPush : io_inputs_1_payload_isPush);
  assign io_output_payload_isPop = (maskRouted_0 ? io_inputs_0_payload_isPop : io_inputs_1_payload_isPop);
  assign io_output_payload_wasWrong = (maskRouted_0 ? io_inputs_0_payload_wasWrong : io_inputs_1_payload_wasWrong);
  assign io_output_payload_badPredictedTarget = (maskRouted_0 ? io_inputs_0_payload_badPredictedTarget : io_inputs_1_payload_badPredictedTarget);
  assign io_output_payload_history = (maskRouted_0 ? io_inputs_0_payload_history : io_inputs_1_payload_history);
  assign io_output_payload_uopId = (maskRouted_0 ? io_inputs_0_payload_uopId : io_inputs_1_payload_uopId);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
    end
  end


endmodule

module StreamArbiter_3 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_op,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [1:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_load,
  input  wire          io_inputs_0_payload_store,
  input  wire          io_inputs_0_payload_atomic,
  input  wire          io_inputs_0_payload_clean,
  input  wire          io_inputs_0_payload_invalidate,
  input  wire [11:0]   io_inputs_0_payload_storeId,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_op,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [1:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_load,
  input  wire          io_inputs_1_payload_store,
  input  wire          io_inputs_1_payload_atomic,
  input  wire          io_inputs_1_payload_clean,
  input  wire          io_inputs_1_payload_invalidate,
  input  wire [11:0]   io_inputs_1_payload_storeId,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_op,
  input  wire [31:0]   io_inputs_2_payload_address,
  input  wire [1:0]    io_inputs_2_payload_size,
  input  wire          io_inputs_2_payload_load,
  input  wire          io_inputs_2_payload_store,
  input  wire          io_inputs_2_payload_atomic,
  input  wire          io_inputs_2_payload_clean,
  input  wire          io_inputs_2_payload_invalidate,
  input  wire [11:0]   io_inputs_2_payload_storeId,
  input  wire          io_inputs_3_valid,
  output wire          io_inputs_3_ready,
  input  wire [2:0]    io_inputs_3_payload_op,
  input  wire [31:0]   io_inputs_3_payload_address,
  input  wire [1:0]    io_inputs_3_payload_size,
  input  wire          io_inputs_3_payload_load,
  input  wire          io_inputs_3_payload_store,
  input  wire          io_inputs_3_payload_atomic,
  input  wire          io_inputs_3_payload_clean,
  input  wire          io_inputs_3_payload_invalidate,
  input  wire [11:0]   io_inputs_3_payload_storeId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_op,
  output wire [31:0]   io_output_payload_address,
  output wire [1:0]    io_output_payload_size,
  output wire          io_output_payload_load,
  output wire          io_output_payload_store,
  output wire          io_output_payload_atomic,
  output wire          io_output_payload_clean,
  output wire          io_output_payload_invalidate,
  output wire [11:0]   io_output_payload_storeId,
  output wire [1:0]    io_chosen,
  output wire [3:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;

  wire       [3:0]    _zz__zz_maskProposal_1_1;
  reg        [2:0]    _zz__zz_io_output_payload_op;
  reg        [31:0]   _zz_io_output_payload_address_3;
  reg        [1:0]    _zz_io_output_payload_size;
  reg                 _zz_io_output_payload_load;
  reg                 _zz_io_output_payload_store;
  reg                 _zz_io_output_payload_atomic;
  reg                 _zz_io_output_payload_clean;
  reg                 _zz_io_output_payload_invalidate;
  reg        [11:0]   _zz_io_output_payload_storeId;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire       [3:0]    _zz_maskProposal_1;
  wire       [3:0]    _zz_maskProposal_1_1;
  wire                _zz_io_output_payload_address;
  wire                _zz_io_output_payload_address_1;
  wire       [1:0]    _zz_io_output_payload_address_2;
  wire       [2:0]    _zz_io_output_payload_op;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;
  `ifndef SYNTHESIS
  reg [95:0] io_inputs_0_payload_op_string;
  reg [95:0] io_inputs_1_payload_op_string;
  reg [95:0] io_inputs_2_payload_op_string;
  reg [95:0] io_inputs_3_payload_op_string;
  reg [95:0] io_output_payload_op_string;
  reg [95:0] _zz_io_output_payload_op_string;
  `endif


  assign _zz__zz_maskProposal_1_1 = (_zz_maskProposal_1 - 4'b0001);
  always @(*) begin
    case(_zz_io_output_payload_address_2)
      2'b00 : begin
        _zz__zz_io_output_payload_op = io_inputs_0_payload_op;
        _zz_io_output_payload_address_3 = io_inputs_0_payload_address;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_load = io_inputs_0_payload_load;
        _zz_io_output_payload_store = io_inputs_0_payload_store;
        _zz_io_output_payload_atomic = io_inputs_0_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_0_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_0_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_0_payload_storeId;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_op = io_inputs_1_payload_op;
        _zz_io_output_payload_address_3 = io_inputs_1_payload_address;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_load = io_inputs_1_payload_load;
        _zz_io_output_payload_store = io_inputs_1_payload_store;
        _zz_io_output_payload_atomic = io_inputs_1_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_1_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_1_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_1_payload_storeId;
      end
      2'b10 : begin
        _zz__zz_io_output_payload_op = io_inputs_2_payload_op;
        _zz_io_output_payload_address_3 = io_inputs_2_payload_address;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_load = io_inputs_2_payload_load;
        _zz_io_output_payload_store = io_inputs_2_payload_store;
        _zz_io_output_payload_atomic = io_inputs_2_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_2_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_2_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_2_payload_storeId;
      end
      default : begin
        _zz__zz_io_output_payload_op = io_inputs_3_payload_op;
        _zz_io_output_payload_address_3 = io_inputs_3_payload_address;
        _zz_io_output_payload_size = io_inputs_3_payload_size;
        _zz_io_output_payload_load = io_inputs_3_payload_load;
        _zz_io_output_payload_store = io_inputs_3_payload_store;
        _zz_io_output_payload_atomic = io_inputs_3_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_3_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_3_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_3_payload_storeId;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_0_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_0_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_0_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_0_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_0_payload_op_string = "PREFETCH    ";
      default : io_inputs_0_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_1_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_1_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_1_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_1_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_1_payload_op_string = "PREFETCH    ";
      default : io_inputs_1_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_2_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_2_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_2_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_2_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_2_payload_op_string = "PREFETCH    ";
      default : io_inputs_2_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_3_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_3_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_3_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_3_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_3_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_3_payload_op_string = "PREFETCH    ";
      default : io_inputs_3_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_op)
      LsuL1CmdOpcode_LSU : io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_output_payload_op_string = "PREFETCH    ";
      default : io_output_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_op)
      LsuL1CmdOpcode_LSU : _zz_io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : _zz_io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : _zz_io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : _zz_io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : _zz_io_output_payload_op_string = "PREFETCH    ";
      default : _zz_io_output_payload_op_string = "????????????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign _zz_maskProposal_1 = {io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}};
  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz__zz_maskProposal_1_1));
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign maskProposal_2 = _zz_maskProposal_1_1[2];
  assign maskProposal_3 = _zz_maskProposal_1_1[3];
  assign io_output_valid = ((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3));
  assign _zz_io_output_payload_address = (maskRouted_1 || maskRouted_3);
  assign _zz_io_output_payload_address_1 = (maskRouted_2 || maskRouted_3);
  assign _zz_io_output_payload_address_2 = {_zz_io_output_payload_address_1,_zz_io_output_payload_address};
  assign _zz_io_output_payload_op = _zz__zz_io_output_payload_op;
  assign io_output_payload_op = _zz_io_output_payload_op;
  assign io_output_payload_address = _zz_io_output_payload_address_3;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_load = _zz_io_output_payload_load;
  assign io_output_payload_store = _zz_io_output_payload_store;
  assign io_output_payload_atomic = _zz_io_output_payload_atomic;
  assign io_output_payload_clean = _zz_io_output_payload_clean;
  assign io_output_payload_invalidate = _zz_io_output_payload_invalidate;
  assign io_output_payload_storeId = _zz_io_output_payload_storeId;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_inputs_2_ready = ((1'b0 || maskRouted_2) && io_output_ready);
  assign io_inputs_3_ready = ((1'b0 || maskRouted_3) && io_output_ready);
  assign io_chosenOH = {maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = (io_chosenOH[1] || _zz_io_chosen);
  assign _zz_io_chosen_2 = (io_chosenOH[2] || _zz_io_chosen);
  assign io_chosen = {_zz_io_chosen_2,_zz_io_chosen_1};
  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
      maskLocked_2 <= maskRouted_2;
      maskLocked_3 <= maskRouted_3;
    end
  end


endmodule

module StreamArbiter_2 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire                io_output_fire;

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskProposal_0 = io_inputs_0_valid;
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
    end
  end


endmodule

module DivRadix (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [63:0]   io_cmd_payload_a,
  input  wire [63:0]   io_cmd_payload_b,
  input  wire          io_cmd_payload_normalized,
  input  wire [4:0]    io_cmd_payload_iterations,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [63:0]   io_rsp_payload_result,
  output wire [63:0]   io_rsp_payload_remain,
  input  wire          clk,
  input  wire          reset
);

  wire       [65:0]   _zz_div3;
  wire       [64:0]   _zz_div3_1;
  wire       [64:0]   _zz_div3_2;
  wire       [15:0]   _zz_shifter_1;
  wire       [31:0]   _zz_shifter_2;
  wire       [47:0]   _zz_shifter_3;
  wire       [61:0]   _zz_shifter_4;
  reg        [4:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix_l45;
  reg        [63:0]   shifter;
  reg        [63:0]   numerator;
  reg        [63:0]   result;
  reg        [65:0]   div1;
  reg        [65:0]   div3;
  wire       [65:0]   div2;
  wire       [65:0]   shifted;
  wire       [66:0]   sub1;
  wire       [66:0]   sub2;
  wire       [66:0]   sub3;
  wire                when_DivRadix_l64;
  reg        [65:0]   _zz_shifter;
  wire                when_DivRadix_l68;
  wire                when_DivRadix_l73;
  wire                when_DivRadix_l77;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  reg                 wasBusy;
  wire                when_DivRadix_l93;

  assign _zz_div3_1 = {1'b0,io_cmd_payload_b};
  assign _zz_div3 = {1'd0, _zz_div3_1};
  assign _zz_div3_2 = ({1'd0,io_cmd_payload_b} <<< 1'd1);
  assign _zz_shifter_1 = io_cmd_payload_a[63 : 48];
  assign _zz_shifter_2 = io_cmd_payload_a[63 : 32];
  assign _zz_shifter_3 = io_cmd_payload_a[63 : 16];
  assign _zz_shifter_4 = io_cmd_payload_a[63 : 2];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix_l45 = (busy && (counter == 5'h1f));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[63 : 62]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign sub2 = ({1'b0,shifted} - {1'b0,div2});
  assign sub3 = ({1'b0,shifted} - {1'b0,div3});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = result;
  assign io_rsp_payload_remain = shifter;
  assign io_cmd_ready = (! busy);
  assign when_DivRadix_l64 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix_l68) begin
      _zz_shifter = sub1[65:0];
    end
    if(when_DivRadix_l73) begin
      _zz_shifter = sub2[65:0];
    end
    if(when_DivRadix_l77) begin
      _zz_shifter = sub3[65:0];
    end
  end

  assign when_DivRadix_l68 = (! sub1[66]);
  assign when_DivRadix_l73 = (! sub2[66]);
  assign when_DivRadix_l77 = (! sub3[66]);
  assign slicesZero_0 = (io_cmd_payload_a[31 : 16] == 16'h0);
  assign slicesZero_1 = (io_cmd_payload_a[47 : 32] == 16'h0);
  assign slicesZero_2 = (io_cmd_payload_a[63 : 48] == 16'h0);
  assign shiftSel = {(&slicesZero_2),{(&{slicesZero_2,slicesZero_1}),(&{slicesZero_2,{slicesZero_1,slicesZero_0}})}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! (|{_zz_sel_2,_zz_sel_1})));
    _zz_sel_4[3] = (_zz_sel[3] && (! (|{_zz_sel_3,{_zz_sel_2,_zz_sel_1}})));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix_l93 = (! busy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      busy <= 1'b0;
      done <= 1'b0;
      wasBusy <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix_l45) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      wasBusy <= busy;
      if(when_DivRadix_l93) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_DivRadix_l64) begin
      counter <= (counter + 5'h01);
      result <= (result <<< 2);
      if(when_DivRadix_l68) begin
        result[1 : 0] <= 2'b01;
      end
      if(when_DivRadix_l73) begin
        result[1 : 0] <= 2'b10;
      end
      if(when_DivRadix_l77) begin
        result[1 : 0] <= 2'b11;
      end
      shifter <= _zz_shifter[63:0];
      numerator <= (numerator <<< 2);
    end
    if(when_DivRadix_l93) begin
      div1 <= {2'd0, io_cmd_payload_b};
      div3 <= (_zz_div3 + {1'b0,_zz_div3_2});
      result <= ((io_cmd_payload_b == 64'h0) ? 64'hffffffffffffffff : 64'h0);
      case(sel)
        2'b11 : begin
          counter <= 5'h0;
          shifter <= 64'h0;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 5'h08;
          shifter <= {48'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        2'b01 : begin
          counter <= 5'h10;
          shifter <= {32'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 32);
        end
        default : begin
          counter <= 5'h18;
          shifter <= {16'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 48);
        end
      endcase
      if(io_cmd_payload_normalized) begin
        counter <= (5'h1f - io_cmd_payload_iterations);
        shifter <= {2'd0, _zz_shifter_4};
        numerator <= (io_cmd_payload_a <<< 62);
      end
    end
  end


endmodule

module StreamArbiter_1 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [51:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [51:0]   io_inputs_1_payload_data,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [51:0]   io_output_payload_data,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire          io_inputs_0_payload_fragment_write,
  input  wire [0:0]    io_inputs_0_payload_fragment_id,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire          io_inputs_1_payload_fragment_write,
  input  wire [0:0]    io_inputs_1_payload_fragment_id,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire          io_output_payload_fragment_write,
  output wire [0:0]    io_output_payload_fragment_id,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                io_output_fire;
  wire                when_Stream_l824;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l824 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_write = (maskRouted_0 ? io_inputs_0_payload_fragment_write : io_inputs_1_payload_fragment_write);
  assign io_output_payload_fragment_id = (maskRouted_0 ? io_inputs_0_payload_fragment_id : io_inputs_1_payload_fragment_id);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l824) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_address,
  input  wire          io_push_payload_unique,
  input  wire [2:0]    io_push_payload_from,
  input  wire [2:0]    io_push_payload_to,
  input  wire [11:0]   io_push_payload_stride,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_address,
  output wire          io_pop_payload_unique,
  output wire [2:0]    io_pop_payload_from,
  output wire [2:0]    io_pop_payload_to,
  output wire [11:0]   io_pop_payload_stride,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire       [50:0]   logic_ram_spinal_port1;
  wire       [50:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_address;
  wire                logic_push_onRam_write_payload_data_unique;
  wire       [2:0]    logic_push_onRam_write_payload_data_from;
  wire       [2:0]    logic_push_onRam_write_payload_data_to;
  wire       [11:0]   logic_push_onRam_write_payload_data_stride;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [31:0]   logic_pop_async_readed_address;
  wire                logic_pop_async_readed_unique;
  wire       [2:0]    logic_pop_async_readed_from;
  wire       [2:0]    logic_pop_async_readed_to;
  wire       [11:0]   logic_pop_async_readed_stride;
  wire       [50:0]   _zz_logic_pop_async_readed_address;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [31:0]   logic_pop_addressGen_translated_payload_address;
  wire                logic_pop_addressGen_translated_payload_unique;
  wire       [2:0]    logic_pop_addressGen_translated_payload_from;
  wire       [2:0]    logic_pop_addressGen_translated_payload_to;
  wire       [11:0]   logic_pop_addressGen_translated_payload_stride;
  (* ram_style = "distributed" *) reg [50:0] logic_ram [0:3];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_stride,{logic_push_onRam_write_payload_data_to,{logic_push_onRam_write_payload_data_from,{logic_push_onRam_write_payload_data_unique,logic_push_onRam_write_payload_data_address}}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data_address = io_push_payload_address;
  assign logic_push_onRam_write_payload_data_unique = io_push_payload_unique;
  assign logic_push_onRam_write_payload_data_from = io_push_payload_from;
  assign logic_push_onRam_write_payload_data_to = io_push_payload_to;
  assign logic_push_onRam_write_payload_data_stride = io_push_payload_stride;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign _zz_logic_pop_async_readed_address = logic_ram_spinal_port1;
  assign logic_pop_async_readed_address = _zz_logic_pop_async_readed_address[31 : 0];
  assign logic_pop_async_readed_unique = _zz_logic_pop_async_readed_address[32];
  assign logic_pop_async_readed_from = _zz_logic_pop_async_readed_address[35 : 33];
  assign logic_pop_async_readed_to = _zz_logic_pop_async_readed_address[38 : 36];
  assign logic_pop_async_readed_stride = _zz_logic_pop_async_readed_address[50 : 39];
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload_address = logic_pop_async_readed_address;
  assign logic_pop_addressGen_translated_payload_unique = logic_pop_async_readed_unique;
  assign logic_pop_addressGen_translated_payload_from = logic_pop_async_readed_from;
  assign logic_pop_addressGen_translated_payload_to = logic_pop_async_readed_to;
  assign logic_pop_addressGen_translated_payload_stride = logic_pop_async_readed_stride;
  assign io_pop_valid = logic_pop_addressGen_translated_valid;
  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  assign io_pop_payload_address = logic_pop_addressGen_translated_payload_address;
  assign io_pop_payload_unique = logic_pop_addressGen_translated_payload_unique;
  assign io_pop_payload_from = logic_pop_addressGen_translated_payload_from;
  assign io_pop_payload_to = logic_pop_addressGen_translated_payload_to;
  assign io_pop_payload_stride = logic_pop_addressGen_translated_payload_stride;
  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
    end
  end


endmodule

module RamSyncMwMux (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [31:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [31:0]   io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [4:0]    io_read_0_cmd_payload,
  output wire [31:0]   io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [4:0]    io_read_1_cmd_payload,
  output wire [31:0]   io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [4:0]    io_read_2_cmd_payload,
  output wire [31:0]   io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [4:0]    io_read_3_cmd_payload,
  output wire [31:0]   io_read_3_rsp,
  input  wire          clk,
  input  wire          reset
);

  reg        [31:0]   ram_0_spinal_port1;
  reg        [31:0]   ram_0_spinal_port2;
  reg        [31:0]   ram_0_spinal_port3;
  reg        [31:0]   ram_0_spinal_port4;
  reg        [31:0]   ram_1_spinal_port1;
  reg        [31:0]   ram_1_spinal_port2;
  reg        [31:0]   ram_1_spinal_port3;
  reg        [31:0]   ram_1_spinal_port4;
  wire       [0:0]    location_io_read_0_rsp;
  wire       [0:0]    location_io_read_1_rsp;
  wire       [0:0]    location_io_read_2_rsp;
  wire       [0:0]    location_io_read_3_rsp;
  reg        [31:0]   _zz_io_read_0_rsp;
  reg        [31:0]   _zz_io_read_1_rsp;
  reg        [31:0]   _zz_io_read_2_rsp;
  reg        [31:0]   _zz_io_read_3_rsp;
  wire       [31:0]   reads_0_reads_0;
  wire       [31:0]   reads_0_reads_1;
  reg        [4:0]    reads_0_addressReg;
  wire       [31:0]   reads_1_reads_0;
  wire       [31:0]   reads_1_reads_1;
  reg        [4:0]    reads_1_addressReg;
  wire       [31:0]   reads_2_reads_0;
  wire       [31:0]   reads_2_reads_1;
  reg        [4:0]    reads_2_addressReg;
  wire       [31:0]   reads_3_reads_0;
  wire       [31:0]   reads_3_reads_1;
  reg        [4:0]    reads_3_addressReg;
  reg [31:0] ram_0 [0:31];
  reg [31:0] ram_1 [0:31];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  always @(posedge clk) begin
    if(io_read_0_cmd_valid) begin
      ram_0_spinal_port1 <= ram_0[io_read_0_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_1_cmd_valid) begin
      ram_0_spinal_port2 <= ram_0[io_read_1_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_2_cmd_valid) begin
      ram_0_spinal_port3 <= ram_0[io_read_2_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_3_cmd_valid) begin
      ram_0_spinal_port4 <= ram_0[io_read_3_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  always @(posedge clk) begin
    if(io_read_0_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[io_read_0_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_1_cmd_valid) begin
      ram_1_spinal_port2 <= ram_1[io_read_1_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_2_cmd_valid) begin
      ram_1_spinal_port3 <= ram_1[io_read_2_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(io_read_3_cmd_valid) begin
      ram_1_spinal_port4 <= ram_1[io_read_3_cmd_payload];
    end
  end

  RamAsyncMwReg location (
    .io_writes_0_valid           (io_writes_0_valid               ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[4:0]), //i
    .io_writes_0_payload_data    (1'b0                            ), //i
    .io_writes_1_valid           (io_writes_1_valid               ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[4:0]), //i
    .io_writes_1_payload_data    (1'b1                            ), //i
    .io_read_0_cmd_valid         (1'b1                            ), //i
    .io_read_0_cmd_payload       (reads_0_addressReg[4:0]         ), //i
    .io_read_0_rsp               (location_io_read_0_rsp          ), //o
    .io_read_1_cmd_valid         (1'b1                            ), //i
    .io_read_1_cmd_payload       (reads_1_addressReg[4:0]         ), //i
    .io_read_1_rsp               (location_io_read_1_rsp          ), //o
    .io_read_2_cmd_valid         (1'b1                            ), //i
    .io_read_2_cmd_payload       (reads_2_addressReg[4:0]         ), //i
    .io_read_2_rsp               (location_io_read_2_rsp          ), //o
    .io_read_3_cmd_valid         (1'b1                            ), //i
    .io_read_3_cmd_payload       (reads_3_addressReg[4:0]         ), //i
    .io_read_3_rsp               (location_io_read_3_rsp          ), //o
    .clk                         (clk                             ), //i
    .reset                       (reset                           )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      1'b0 : _zz_io_read_0_rsp = reads_0_reads_0;
      default : _zz_io_read_0_rsp = reads_0_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_1_rsp)
      1'b0 : _zz_io_read_1_rsp = reads_1_reads_0;
      default : _zz_io_read_1_rsp = reads_1_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_2_rsp)
      1'b0 : _zz_io_read_2_rsp = reads_2_reads_0;
      default : _zz_io_read_2_rsp = reads_2_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_3_rsp)
      1'b0 : _zz_io_read_3_rsp = reads_3_reads_0;
      default : _zz_io_read_3_rsp = reads_3_reads_1;
    endcase
  end

  assign reads_0_reads_0 = ram_0_spinal_port1;
  assign reads_0_reads_1 = ram_1_spinal_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign reads_1_reads_0 = ram_0_spinal_port2;
  assign reads_1_reads_1 = ram_1_spinal_port2;
  assign io_read_1_rsp = _zz_io_read_1_rsp;
  assign reads_2_reads_0 = ram_0_spinal_port3;
  assign reads_2_reads_1 = ram_1_spinal_port3;
  assign io_read_2_rsp = _zz_io_read_2_rsp;
  assign reads_3_reads_0 = ram_0_spinal_port4;
  assign reads_3_reads_1 = ram_1_spinal_port4;
  assign io_read_3_rsp = _zz_io_read_3_rsp;
  always @(posedge clk) begin
    if(io_read_0_cmd_valid) begin
      reads_0_addressReg <= io_read_0_cmd_payload;
    end
    if(io_read_1_cmd_valid) begin
      reads_1_addressReg <= io_read_1_cmd_payload;
    end
    if(io_read_2_cmd_valid) begin
      reads_2_addressReg <= io_read_2_cmd_payload;
    end
    if(io_read_3_cmd_valid) begin
      reads_3_addressReg <= io_read_3_cmd_payload;
    end
  end


endmodule

module RamAsyncMwReg (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [4:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [4:0]    io_read_1_cmd_payload,
  output wire [0:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [4:0]    io_read_2_cmd_payload,
  output wire [0:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [4:0]    io_read_3_cmd_payload,
  output wire [0:0]    io_read_3_rsp,
  input  wire          clk,
  input  wire          reset
);

  reg        [0:0]    _zz_io_read_0_rsp;
  reg        [0:0]    _zz_io_read_1_rsp;
  reg        [0:0]    _zz_io_read_2_rsp;
  reg        [0:0]    _zz_io_read_3_rsp;
  reg        [0:0]    ram_0;
  reg        [0:0]    ram_1;
  reg        [0:0]    ram_2;
  reg        [0:0]    ram_3;
  reg        [0:0]    ram_4;
  reg        [0:0]    ram_5;
  reg        [0:0]    ram_6;
  reg        [0:0]    ram_7;
  reg        [0:0]    ram_8;
  reg        [0:0]    ram_9;
  reg        [0:0]    ram_10;
  reg        [0:0]    ram_11;
  reg        [0:0]    ram_12;
  reg        [0:0]    ram_13;
  reg        [0:0]    ram_14;
  reg        [0:0]    ram_15;
  reg        [0:0]    ram_16;
  reg        [0:0]    ram_17;
  reg        [0:0]    ram_18;
  reg        [0:0]    ram_19;
  reg        [0:0]    ram_20;
  reg        [0:0]    ram_21;
  reg        [0:0]    ram_22;
  reg        [0:0]    ram_23;
  reg        [0:0]    ram_24;
  reg        [0:0]    ram_25;
  reg        [0:0]    ram_26;
  reg        [0:0]    ram_27;
  reg        [0:0]    ram_28;
  reg        [0:0]    ram_29;
  reg        [0:0]    ram_30;
  reg        [0:0]    ram_31;
  wire       [31:0]   _zz_1;
  wire       [0:0]    _zz_ram_0;
  wire       [31:0]   _zz_2;
  wire       [0:0]    _zz_ram_0_1;

  initial begin
  `ifndef SYNTHESIS
    ram_0 = {$urandom};
    ram_1 = {$urandom};
    ram_2 = {$urandom};
    ram_3 = {$urandom};
    ram_4 = {$urandom};
    ram_5 = {$urandom};
    ram_6 = {$urandom};
    ram_7 = {$urandom};
    ram_8 = {$urandom};
    ram_9 = {$urandom};
    ram_10 = {$urandom};
    ram_11 = {$urandom};
    ram_12 = {$urandom};
    ram_13 = {$urandom};
    ram_14 = {$urandom};
    ram_15 = {$urandom};
    ram_16 = {$urandom};
    ram_17 = {$urandom};
    ram_18 = {$urandom};
    ram_19 = {$urandom};
    ram_20 = {$urandom};
    ram_21 = {$urandom};
    ram_22 = {$urandom};
    ram_23 = {$urandom};
    ram_24 = {$urandom};
    ram_25 = {$urandom};
    ram_26 = {$urandom};
    ram_27 = {$urandom};
    ram_28 = {$urandom};
    ram_29 = {$urandom};
    ram_30 = {$urandom};
    ram_31 = {$urandom};
  `endif
  end

  always @(*) begin
    case(io_read_0_cmd_payload)
      5'b00000 : _zz_io_read_0_rsp = ram_0;
      5'b00001 : _zz_io_read_0_rsp = ram_1;
      5'b00010 : _zz_io_read_0_rsp = ram_2;
      5'b00011 : _zz_io_read_0_rsp = ram_3;
      5'b00100 : _zz_io_read_0_rsp = ram_4;
      5'b00101 : _zz_io_read_0_rsp = ram_5;
      5'b00110 : _zz_io_read_0_rsp = ram_6;
      5'b00111 : _zz_io_read_0_rsp = ram_7;
      5'b01000 : _zz_io_read_0_rsp = ram_8;
      5'b01001 : _zz_io_read_0_rsp = ram_9;
      5'b01010 : _zz_io_read_0_rsp = ram_10;
      5'b01011 : _zz_io_read_0_rsp = ram_11;
      5'b01100 : _zz_io_read_0_rsp = ram_12;
      5'b01101 : _zz_io_read_0_rsp = ram_13;
      5'b01110 : _zz_io_read_0_rsp = ram_14;
      5'b01111 : _zz_io_read_0_rsp = ram_15;
      5'b10000 : _zz_io_read_0_rsp = ram_16;
      5'b10001 : _zz_io_read_0_rsp = ram_17;
      5'b10010 : _zz_io_read_0_rsp = ram_18;
      5'b10011 : _zz_io_read_0_rsp = ram_19;
      5'b10100 : _zz_io_read_0_rsp = ram_20;
      5'b10101 : _zz_io_read_0_rsp = ram_21;
      5'b10110 : _zz_io_read_0_rsp = ram_22;
      5'b10111 : _zz_io_read_0_rsp = ram_23;
      5'b11000 : _zz_io_read_0_rsp = ram_24;
      5'b11001 : _zz_io_read_0_rsp = ram_25;
      5'b11010 : _zz_io_read_0_rsp = ram_26;
      5'b11011 : _zz_io_read_0_rsp = ram_27;
      5'b11100 : _zz_io_read_0_rsp = ram_28;
      5'b11101 : _zz_io_read_0_rsp = ram_29;
      5'b11110 : _zz_io_read_0_rsp = ram_30;
      default : _zz_io_read_0_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_1_cmd_payload)
      5'b00000 : _zz_io_read_1_rsp = ram_0;
      5'b00001 : _zz_io_read_1_rsp = ram_1;
      5'b00010 : _zz_io_read_1_rsp = ram_2;
      5'b00011 : _zz_io_read_1_rsp = ram_3;
      5'b00100 : _zz_io_read_1_rsp = ram_4;
      5'b00101 : _zz_io_read_1_rsp = ram_5;
      5'b00110 : _zz_io_read_1_rsp = ram_6;
      5'b00111 : _zz_io_read_1_rsp = ram_7;
      5'b01000 : _zz_io_read_1_rsp = ram_8;
      5'b01001 : _zz_io_read_1_rsp = ram_9;
      5'b01010 : _zz_io_read_1_rsp = ram_10;
      5'b01011 : _zz_io_read_1_rsp = ram_11;
      5'b01100 : _zz_io_read_1_rsp = ram_12;
      5'b01101 : _zz_io_read_1_rsp = ram_13;
      5'b01110 : _zz_io_read_1_rsp = ram_14;
      5'b01111 : _zz_io_read_1_rsp = ram_15;
      5'b10000 : _zz_io_read_1_rsp = ram_16;
      5'b10001 : _zz_io_read_1_rsp = ram_17;
      5'b10010 : _zz_io_read_1_rsp = ram_18;
      5'b10011 : _zz_io_read_1_rsp = ram_19;
      5'b10100 : _zz_io_read_1_rsp = ram_20;
      5'b10101 : _zz_io_read_1_rsp = ram_21;
      5'b10110 : _zz_io_read_1_rsp = ram_22;
      5'b10111 : _zz_io_read_1_rsp = ram_23;
      5'b11000 : _zz_io_read_1_rsp = ram_24;
      5'b11001 : _zz_io_read_1_rsp = ram_25;
      5'b11010 : _zz_io_read_1_rsp = ram_26;
      5'b11011 : _zz_io_read_1_rsp = ram_27;
      5'b11100 : _zz_io_read_1_rsp = ram_28;
      5'b11101 : _zz_io_read_1_rsp = ram_29;
      5'b11110 : _zz_io_read_1_rsp = ram_30;
      default : _zz_io_read_1_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_2_cmd_payload)
      5'b00000 : _zz_io_read_2_rsp = ram_0;
      5'b00001 : _zz_io_read_2_rsp = ram_1;
      5'b00010 : _zz_io_read_2_rsp = ram_2;
      5'b00011 : _zz_io_read_2_rsp = ram_3;
      5'b00100 : _zz_io_read_2_rsp = ram_4;
      5'b00101 : _zz_io_read_2_rsp = ram_5;
      5'b00110 : _zz_io_read_2_rsp = ram_6;
      5'b00111 : _zz_io_read_2_rsp = ram_7;
      5'b01000 : _zz_io_read_2_rsp = ram_8;
      5'b01001 : _zz_io_read_2_rsp = ram_9;
      5'b01010 : _zz_io_read_2_rsp = ram_10;
      5'b01011 : _zz_io_read_2_rsp = ram_11;
      5'b01100 : _zz_io_read_2_rsp = ram_12;
      5'b01101 : _zz_io_read_2_rsp = ram_13;
      5'b01110 : _zz_io_read_2_rsp = ram_14;
      5'b01111 : _zz_io_read_2_rsp = ram_15;
      5'b10000 : _zz_io_read_2_rsp = ram_16;
      5'b10001 : _zz_io_read_2_rsp = ram_17;
      5'b10010 : _zz_io_read_2_rsp = ram_18;
      5'b10011 : _zz_io_read_2_rsp = ram_19;
      5'b10100 : _zz_io_read_2_rsp = ram_20;
      5'b10101 : _zz_io_read_2_rsp = ram_21;
      5'b10110 : _zz_io_read_2_rsp = ram_22;
      5'b10111 : _zz_io_read_2_rsp = ram_23;
      5'b11000 : _zz_io_read_2_rsp = ram_24;
      5'b11001 : _zz_io_read_2_rsp = ram_25;
      5'b11010 : _zz_io_read_2_rsp = ram_26;
      5'b11011 : _zz_io_read_2_rsp = ram_27;
      5'b11100 : _zz_io_read_2_rsp = ram_28;
      5'b11101 : _zz_io_read_2_rsp = ram_29;
      5'b11110 : _zz_io_read_2_rsp = ram_30;
      default : _zz_io_read_2_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_3_cmd_payload)
      5'b00000 : _zz_io_read_3_rsp = ram_0;
      5'b00001 : _zz_io_read_3_rsp = ram_1;
      5'b00010 : _zz_io_read_3_rsp = ram_2;
      5'b00011 : _zz_io_read_3_rsp = ram_3;
      5'b00100 : _zz_io_read_3_rsp = ram_4;
      5'b00101 : _zz_io_read_3_rsp = ram_5;
      5'b00110 : _zz_io_read_3_rsp = ram_6;
      5'b00111 : _zz_io_read_3_rsp = ram_7;
      5'b01000 : _zz_io_read_3_rsp = ram_8;
      5'b01001 : _zz_io_read_3_rsp = ram_9;
      5'b01010 : _zz_io_read_3_rsp = ram_10;
      5'b01011 : _zz_io_read_3_rsp = ram_11;
      5'b01100 : _zz_io_read_3_rsp = ram_12;
      5'b01101 : _zz_io_read_3_rsp = ram_13;
      5'b01110 : _zz_io_read_3_rsp = ram_14;
      5'b01111 : _zz_io_read_3_rsp = ram_15;
      5'b10000 : _zz_io_read_3_rsp = ram_16;
      5'b10001 : _zz_io_read_3_rsp = ram_17;
      5'b10010 : _zz_io_read_3_rsp = ram_18;
      5'b10011 : _zz_io_read_3_rsp = ram_19;
      5'b10100 : _zz_io_read_3_rsp = ram_20;
      5'b10101 : _zz_io_read_3_rsp = ram_21;
      5'b10110 : _zz_io_read_3_rsp = ram_22;
      5'b10111 : _zz_io_read_3_rsp = ram_23;
      5'b11000 : _zz_io_read_3_rsp = ram_24;
      5'b11001 : _zz_io_read_3_rsp = ram_25;
      5'b11010 : _zz_io_read_3_rsp = ram_26;
      5'b11011 : _zz_io_read_3_rsp = ram_27;
      5'b11100 : _zz_io_read_3_rsp = ram_28;
      5'b11101 : _zz_io_read_3_rsp = ram_29;
      5'b11110 : _zz_io_read_3_rsp = ram_30;
      default : _zz_io_read_3_rsp = ram_31;
    endcase
  end

  assign _zz_1 = ({31'd0,1'b1} <<< io_writes_0_payload_address);
  assign _zz_ram_0 = io_writes_0_payload_data;
  assign _zz_2 = ({31'd0,1'b1} <<< io_writes_1_payload_address);
  assign _zz_ram_0_1 = io_writes_1_payload_data;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign io_read_1_rsp = _zz_io_read_1_rsp;
  assign io_read_2_rsp = _zz_io_read_2_rsp;
  assign io_read_3_rsp = _zz_io_read_3_rsp;
  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      if(_zz_1[0]) begin
        ram_0 <= _zz_ram_0;
      end
      if(_zz_1[1]) begin
        ram_1 <= _zz_ram_0;
      end
      if(_zz_1[2]) begin
        ram_2 <= _zz_ram_0;
      end
      if(_zz_1[3]) begin
        ram_3 <= _zz_ram_0;
      end
      if(_zz_1[4]) begin
        ram_4 <= _zz_ram_0;
      end
      if(_zz_1[5]) begin
        ram_5 <= _zz_ram_0;
      end
      if(_zz_1[6]) begin
        ram_6 <= _zz_ram_0;
      end
      if(_zz_1[7]) begin
        ram_7 <= _zz_ram_0;
      end
      if(_zz_1[8]) begin
        ram_8 <= _zz_ram_0;
      end
      if(_zz_1[9]) begin
        ram_9 <= _zz_ram_0;
      end
      if(_zz_1[10]) begin
        ram_10 <= _zz_ram_0;
      end
      if(_zz_1[11]) begin
        ram_11 <= _zz_ram_0;
      end
      if(_zz_1[12]) begin
        ram_12 <= _zz_ram_0;
      end
      if(_zz_1[13]) begin
        ram_13 <= _zz_ram_0;
      end
      if(_zz_1[14]) begin
        ram_14 <= _zz_ram_0;
      end
      if(_zz_1[15]) begin
        ram_15 <= _zz_ram_0;
      end
      if(_zz_1[16]) begin
        ram_16 <= _zz_ram_0;
      end
      if(_zz_1[17]) begin
        ram_17 <= _zz_ram_0;
      end
      if(_zz_1[18]) begin
        ram_18 <= _zz_ram_0;
      end
      if(_zz_1[19]) begin
        ram_19 <= _zz_ram_0;
      end
      if(_zz_1[20]) begin
        ram_20 <= _zz_ram_0;
      end
      if(_zz_1[21]) begin
        ram_21 <= _zz_ram_0;
      end
      if(_zz_1[22]) begin
        ram_22 <= _zz_ram_0;
      end
      if(_zz_1[23]) begin
        ram_23 <= _zz_ram_0;
      end
      if(_zz_1[24]) begin
        ram_24 <= _zz_ram_0;
      end
      if(_zz_1[25]) begin
        ram_25 <= _zz_ram_0;
      end
      if(_zz_1[26]) begin
        ram_26 <= _zz_ram_0;
      end
      if(_zz_1[27]) begin
        ram_27 <= _zz_ram_0;
      end
      if(_zz_1[28]) begin
        ram_28 <= _zz_ram_0;
      end
      if(_zz_1[29]) begin
        ram_29 <= _zz_ram_0;
      end
      if(_zz_1[30]) begin
        ram_30 <= _zz_ram_0;
      end
      if(_zz_1[31]) begin
        ram_31 <= _zz_ram_0;
      end
    end
    if(io_writes_1_valid) begin
      if(_zz_2[0]) begin
        ram_0 <= _zz_ram_0_1;
      end
      if(_zz_2[1]) begin
        ram_1 <= _zz_ram_0_1;
      end
      if(_zz_2[2]) begin
        ram_2 <= _zz_ram_0_1;
      end
      if(_zz_2[3]) begin
        ram_3 <= _zz_ram_0_1;
      end
      if(_zz_2[4]) begin
        ram_4 <= _zz_ram_0_1;
      end
      if(_zz_2[5]) begin
        ram_5 <= _zz_ram_0_1;
      end
      if(_zz_2[6]) begin
        ram_6 <= _zz_ram_0_1;
      end
      if(_zz_2[7]) begin
        ram_7 <= _zz_ram_0_1;
      end
      if(_zz_2[8]) begin
        ram_8 <= _zz_ram_0_1;
      end
      if(_zz_2[9]) begin
        ram_9 <= _zz_ram_0_1;
      end
      if(_zz_2[10]) begin
        ram_10 <= _zz_ram_0_1;
      end
      if(_zz_2[11]) begin
        ram_11 <= _zz_ram_0_1;
      end
      if(_zz_2[12]) begin
        ram_12 <= _zz_ram_0_1;
      end
      if(_zz_2[13]) begin
        ram_13 <= _zz_ram_0_1;
      end
      if(_zz_2[14]) begin
        ram_14 <= _zz_ram_0_1;
      end
      if(_zz_2[15]) begin
        ram_15 <= _zz_ram_0_1;
      end
      if(_zz_2[16]) begin
        ram_16 <= _zz_ram_0_1;
      end
      if(_zz_2[17]) begin
        ram_17 <= _zz_ram_0_1;
      end
      if(_zz_2[18]) begin
        ram_18 <= _zz_ram_0_1;
      end
      if(_zz_2[19]) begin
        ram_19 <= _zz_ram_0_1;
      end
      if(_zz_2[20]) begin
        ram_20 <= _zz_ram_0_1;
      end
      if(_zz_2[21]) begin
        ram_21 <= _zz_ram_0_1;
      end
      if(_zz_2[22]) begin
        ram_22 <= _zz_ram_0_1;
      end
      if(_zz_2[23]) begin
        ram_23 <= _zz_ram_0_1;
      end
      if(_zz_2[24]) begin
        ram_24 <= _zz_ram_0_1;
      end
      if(_zz_2[25]) begin
        ram_25 <= _zz_ram_0_1;
      end
      if(_zz_2[26]) begin
        ram_26 <= _zz_ram_0_1;
      end
      if(_zz_2[27]) begin
        ram_27 <= _zz_ram_0_1;
      end
      if(_zz_2[28]) begin
        ram_28 <= _zz_ram_0_1;
      end
      if(_zz_2[29]) begin
        ram_29 <= _zz_ram_0_1;
      end
      if(_zz_2[30]) begin
        ram_30 <= _zz_ram_0_1;
      end
      if(_zz_2[31]) begin
        ram_31 <= _zz_ram_0_1;
      end
    end
  end


endmodule
